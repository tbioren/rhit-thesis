module individual (
    (* keep *) input in0, in1, in2, in3, in4, in5, in6, in7, in8, in9,
    (* keep *) output out0, out1, out2, out3, out4, out5, out6, out7, out8, out9);
    wire x1_y1;
    wire x2_y1;
    wire x3_y1;
    wire x4_y1;
    wire x5_y1;
    wire x7_y1;
    wire x8_y1;
    wire x9_y1;
    wire x10_y1;
    wire x11_y1;
    wire x1_y2;
    wire x2_y2;
    wire x3_y2;
    wire x4_y2;
    wire x5_y2;
    wire x7_y2;
    wire x8_y2;
    wire x9_y2;
    wire x10_y2;
    wire x11_y2;
    wire x1_y3;
    wire x2_y3;
    wire x3_y3;
    wire x4_y3;
    wire x5_y3;
    wire x7_y3;
    wire x8_y3;
    wire x9_y3;
    wire x10_y3;
    wire x11_y3;
    wire x1_y4;
    wire x2_y4;
    wire x3_y4;
    wire x4_y4;
    wire x5_y4;
    wire x7_y4;
    wire x8_y4;
    wire x9_y4;
    wire x10_y4;
    wire x11_y4;
    wire x1_y5;
    wire x2_y5;
    wire x3_y5;
    wire x4_y5;
    wire x5_y5;
    wire x7_y5;
    wire x8_y5;
    wire x9_y5;
    wire x10_y5;
    wire x11_y5;
    wire x1_y6;
    wire x2_y6;
    wire x3_y6;
    wire x4_y6;
    wire x5_y6;
    wire x7_y6;
    wire x8_y6;
    wire x9_y6;
    wire x10_y6;
    wire x11_y6;
    wire x1_y7;
    wire x2_y7;
    wire x3_y7;
    wire x4_y7;
    wire x5_y7;
    wire x7_y7;
    wire x8_y7;
    wire x9_y7;
    wire x10_y7;
    wire x11_y7;
    wire x1_y8;
    wire x2_y8;
    wire x3_y8;
    wire x4_y8;
    wire x5_y8;
    wire x7_y8;
    wire x8_y8;
    wire x9_y8;
    wire x10_y8;
    wire x11_y8;
    wire x1_y9;
    wire x2_y9;
    wire x3_y9;
    wire x4_y9;
    wire x5_y9;
    wire x7_y9;
    wire x8_y9;
    wire x9_y9;
    wire x10_y9;
    wire x11_y9;
    wire x1_y10;
    wire x2_y10;
    wire x3_y10;
    wire x4_y10;
    wire x5_y10;
    wire x7_y10;
    wire x8_y10;
    wire x9_y10;
    wire x10_y10;
    wire x11_y10;

    (* keep, dont_touch *)
    (* BEL = "X1/Y1/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000007)
    ) lut_1_1 (
        .O(x1_y1),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X2/Y1/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000008)
    ) lut_2_1 (
        .O(x2_y1),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X3/Y1/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000008)
    ) lut_3_1 (
        .O(x3_y1),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X4/Y1/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000007)
    ) lut_4_1 (
        .O(x4_y1),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X5/Y1/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000015)
    ) lut_5_1 (
        .O(x5_y1),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X7/Y1/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000005)
    ) lut_7_1 (
        .O(x7_y1),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X8/Y1/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000009)
    ) lut_8_1 (
        .O(x8_y1),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X9/Y1/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000001)
    ) lut_9_1 (
        .O(x9_y1),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X10/Y1/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000015)
    ) lut_10_1 (
        .O(x10_y1),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X11/Y1/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000001)
    ) lut_11_1 (
        .O(x11_y1),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X1/Y1/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000009)
    ) lut_1_2 (
        .O(x1_y2),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X2/Y1/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000002)
    ) lut_2_2 (
        .O(x2_y2),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X3/Y1/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000010)
    ) lut_3_2 (
        .O(x3_y2),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X4/Y1/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000005)
    ) lut_4_2 (
        .O(x4_y2),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X5/Y1/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000010)
    ) lut_5_2 (
        .O(x5_y2),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X7/Y1/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000006)
    ) lut_7_2 (
        .O(x7_y2),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X8/Y1/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000003)
    ) lut_8_2 (
        .O(x8_y2),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X9/Y1/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000003)
    ) lut_9_2 (
        .O(x9_y2),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X10/Y1/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000012)
    ) lut_10_2 (
        .O(x10_y2),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X11/Y1/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000014)
    ) lut_11_2 (
        .O(x11_y2),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X1/Y1/lc2" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000013)
    ) lut_1_3 (
        .O(x1_y3),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X2/Y1/lc2" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000014)
    ) lut_2_3 (
        .O(x2_y3),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X3/Y1/lc2" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000009)
    ) lut_3_3 (
        .O(x3_y3),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X4/Y1/lc2" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000010)
    ) lut_4_3 (
        .O(x4_y3),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X5/Y1/lc2" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000004)
    ) lut_5_3 (
        .O(x5_y3),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X7/Y1/lc2" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000000)
    ) lut_7_3 (
        .O(x7_y3),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X8/Y1/lc2" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000006)
    ) lut_8_3 (
        .O(x8_y3),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X9/Y1/lc2" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000013)
    ) lut_9_3 (
        .O(x9_y3),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X10/Y1/lc2" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000014)
    ) lut_10_3 (
        .O(x10_y3),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X11/Y1/lc2" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000014)
    ) lut_11_3 (
        .O(x11_y3),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X1/Y1/lc3" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000004)
    ) lut_1_4 (
        .O(x1_y4),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X2/Y1/lc3" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000007)
    ) lut_2_4 (
        .O(x2_y4),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X3/Y1/lc3" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000011)
    ) lut_3_4 (
        .O(x3_y4),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X4/Y1/lc3" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000006)
    ) lut_4_4 (
        .O(x4_y4),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X5/Y1/lc3" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000010)
    ) lut_5_4 (
        .O(x5_y4),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X7/Y1/lc3" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000006)
    ) lut_7_4 (
        .O(x7_y4),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X8/Y1/lc3" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000009)
    ) lut_8_4 (
        .O(x8_y4),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X9/Y1/lc3" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000001)
    ) lut_9_4 (
        .O(x9_y4),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X10/Y1/lc3" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000000)
    ) lut_10_4 (
        .O(x10_y4),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X11/Y1/lc3" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000014)
    ) lut_11_4 (
        .O(x11_y4),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X1/Y1/lc4" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000012)
    ) lut_1_5 (
        .O(x1_y5),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X2/Y1/lc4" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000007)
    ) lut_2_5 (
        .O(x2_y5),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X3/Y1/lc4" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000001)
    ) lut_3_5 (
        .O(x3_y5),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X4/Y1/lc4" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000003)
    ) lut_4_5 (
        .O(x4_y5),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X5/Y1/lc4" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000007)
    ) lut_5_5 (
        .O(x5_y5),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X7/Y1/lc4" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000015)
    ) lut_7_5 (
        .O(x7_y5),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X8/Y1/lc4" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000008)
    ) lut_8_5 (
        .O(x8_y5),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X9/Y1/lc4" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000013)
    ) lut_9_5 (
        .O(x9_y5),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X10/Y1/lc4" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000000)
    ) lut_10_5 (
        .O(x10_y5),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X11/Y1/lc4" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000014)
    ) lut_11_5 (
        .O(x11_y5),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X1/Y1/lc5" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000004)
    ) lut_1_6 (
        .O(x1_y6),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X2/Y1/lc5" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000001)
    ) lut_2_6 (
        .O(x2_y6),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X3/Y1/lc5" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000011)
    ) lut_3_6 (
        .O(x3_y6),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X4/Y1/lc5" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000007)
    ) lut_4_6 (
        .O(x4_y6),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X5/Y1/lc5" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000005)
    ) lut_5_6 (
        .O(x5_y6),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X7/Y1/lc5" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000005)
    ) lut_7_6 (
        .O(x7_y6),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X8/Y1/lc5" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000008)
    ) lut_8_6 (
        .O(x8_y6),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X9/Y1/lc5" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000013)
    ) lut_9_6 (
        .O(x9_y6),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X10/Y1/lc5" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000001)
    ) lut_10_6 (
        .O(x10_y6),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X11/Y1/lc5" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000015)
    ) lut_11_6 (
        .O(x11_y6),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X1/Y1/lc6" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000005)
    ) lut_1_7 (
        .O(x1_y7),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X2/Y1/lc6" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000012)
    ) lut_2_7 (
        .O(x2_y7),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X3/Y1/lc6" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000011)
    ) lut_3_7 (
        .O(x3_y7),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X4/Y1/lc6" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000010)
    ) lut_4_7 (
        .O(x4_y7),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X5/Y1/lc6" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000003)
    ) lut_5_7 (
        .O(x5_y7),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X7/Y1/lc6" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000010)
    ) lut_7_7 (
        .O(x7_y7),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X8/Y1/lc6" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000013)
    ) lut_8_7 (
        .O(x8_y7),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X9/Y1/lc6" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000000)
    ) lut_9_7 (
        .O(x9_y7),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X10/Y1/lc6" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000008)
    ) lut_10_7 (
        .O(x10_y7),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X11/Y1/lc6" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000006)
    ) lut_11_7 (
        .O(x11_y7),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X1/Y1/lc7" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000009)
    ) lut_1_8 (
        .O(x1_y8),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X2/Y1/lc7" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000002)
    ) lut_2_8 (
        .O(x2_y8),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X3/Y1/lc7" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000003)
    ) lut_3_8 (
        .O(x3_y8),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X4/Y1/lc7" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000007)
    ) lut_4_8 (
        .O(x4_y8),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X5/Y1/lc7" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000009)
    ) lut_5_8 (
        .O(x5_y8),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X7/Y1/lc7" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000003)
    ) lut_7_8 (
        .O(x7_y8),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X8/Y1/lc7" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000013)
    ) lut_8_8 (
        .O(x8_y8),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X9/Y1/lc7" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000015)
    ) lut_9_8 (
        .O(x9_y8),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X10/Y1/lc7" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000005)
    ) lut_10_8 (
        .O(x10_y8),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X11/Y1/lc7" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000014)
    ) lut_11_8 (
        .O(x11_y8),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X1/Y2/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000013)
    ) lut_1_9 (
        .O(x1_y9),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X2/Y2/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000007)
    ) lut_2_9 (
        .O(x2_y9),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X3/Y2/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000002)
    ) lut_3_9 (
        .O(x3_y9),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X4/Y2/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000011)
    ) lut_4_9 (
        .O(x4_y9),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X5/Y2/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000004)
    ) lut_5_9 (
        .O(x5_y9),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X7/Y2/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000008)
    ) lut_7_9 (
        .O(x7_y9),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X8/Y2/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000015)
    ) lut_8_9 (
        .O(x8_y9),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X9/Y2/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000010)
    ) lut_9_9 (
        .O(x9_y9),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X10/Y2/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000012)
    ) lut_10_9 (
        .O(x10_y9),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X11/Y2/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000014)
    ) lut_11_9 (
        .O(x11_y9),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X1/Y2/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000010)
    ) lut_1_10 (
        .O(x1_y10),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X2/Y2/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000013)
    ) lut_2_10 (
        .O(x2_y10),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X3/Y2/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000011)
    ) lut_3_10 (
        .O(x3_y10),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X4/Y2/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000007)
    ) lut_4_10 (
        .O(x4_y10),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X5/Y2/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000001)
    ) lut_5_10 (
        .O(x5_y10),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X7/Y2/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000006)
    ) lut_7_10 (
        .O(x7_y10),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X8/Y2/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000007)
    ) lut_8_10 (
        .O(x8_y10),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X9/Y2/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000013)
    ) lut_9_10 (
        .O(x9_y10),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X10/Y2/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000010)
    ) lut_10_10 (
        .O(x10_y10),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X11/Y2/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000003)
    ) lut_11_10 (
        .O(x11_y10),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
endmodule
