module cgp_module (
    (* keep *) input in0, in1, in2, in3, in4, in5, in6, in7, in8, in9,
    (* keep *) output out0, out1, out2, out3, out4, out5, out6, out7, out8, out9);

    (* keep *) wire x0_y0, x1_y0, x2_y0, x3_y0, x4_y0, x5_y0, x6_y0, x7_y0, x8_y0, x9_y0, x10_y0, x11_y0, x12_y0, x13_y0, x14_y0, x15_y0, x16_y0, x17_y0, x18_y0, x19_y0, x20_y0, x21_y0, x22_y0, x23_y0, x24_y0, x25_y0, x26_y0, x27_y0, x28_y0, x29_y0, x30_y0, x31_y0, x32_y0, x33_y0, x34_y0, x35_y0, x36_y0, x37_y0, x38_y0, x39_y0, x40_y0, x41_y0, x42_y0, x43_y0, x44_y0, x45_y0, x46_y0, x47_y0, x48_y0, x49_y0, x50_y0, x51_y0, x52_y0, x53_y0, x54_y0, x55_y0, x56_y0, x57_y0, x58_y0, x59_y0, x60_y0, x61_y0, x0_y1, x1_y1, x2_y1, x3_y1, x4_y1, x5_y1, x6_y1, x7_y1, x8_y1, x9_y1, x10_y1, x11_y1, x12_y1, x13_y1, x14_y1, x15_y1, x16_y1, x17_y1, x18_y1, x19_y1, x20_y1, x21_y1, x22_y1, x23_y1, x24_y1, x25_y1, x26_y1, x27_y1, x28_y1, x29_y1, x30_y1, x31_y1, x32_y1, x33_y1, x34_y1, x35_y1, x36_y1, x37_y1, x38_y1, x39_y1, x40_y1, x41_y1, x42_y1, x43_y1, x44_y1, x45_y1, x46_y1, x47_y1, x48_y1, x49_y1, x50_y1, x51_y1, x52_y1, x53_y1, x54_y1, x55_y1, x56_y1, x57_y1, x58_y1, x59_y1, x60_y1, x61_y1, x0_y2, x1_y2, x2_y2, x3_y2, x4_y2, x5_y2, x6_y2, x7_y2, x8_y2, x9_y2, x10_y2, x11_y2, x12_y2, x13_y2, x14_y2, x15_y2, x16_y2, x17_y2, x18_y2, x19_y2, x20_y2, x21_y2, x22_y2, x23_y2, x24_y2, x25_y2, x26_y2, x27_y2, x28_y2, x29_y2, x30_y2, x31_y2, x32_y2, x33_y2, x34_y2, x35_y2, x36_y2, x37_y2, x38_y2, x39_y2, x40_y2, x41_y2, x42_y2, x43_y2, x44_y2, x45_y2, x46_y2, x47_y2, x48_y2, x49_y2, x50_y2, x51_y2, x52_y2, x53_y2, x54_y2, x55_y2, x56_y2, x57_y2, x58_y2, x59_y2, x60_y2, x61_y2, x0_y3, x1_y3, x2_y3, x3_y3, x4_y3, x5_y3, x6_y3, x7_y3, x8_y3, x9_y3, x10_y3, x11_y3, x12_y3, x13_y3, x14_y3, x15_y3, x16_y3, x17_y3, x18_y3, x19_y3, x20_y3, x21_y3, x22_y3, x23_y3, x24_y3, x25_y3, x26_y3, x27_y3, x28_y3, x29_y3, x30_y3, x31_y3, x32_y3, x33_y3, x34_y3, x35_y3, x36_y3, x37_y3, x38_y3, x39_y3, x40_y3, x41_y3, x42_y3, x43_y3, x44_y3, x45_y3, x46_y3, x47_y3, x48_y3, x49_y3, x50_y3, x51_y3, x52_y3, x53_y3, x54_y3, x55_y3, x56_y3, x57_y3, x58_y3, x59_y3, x60_y3, x61_y3, x0_y4, x1_y4, x2_y4, x3_y4, x4_y4, x5_y4, x6_y4, x7_y4, x8_y4, x9_y4, x10_y4, x11_y4, x12_y4, x13_y4, x14_y4, x15_y4, x16_y4, x17_y4, x18_y4, x19_y4, x20_y4, x21_y4, x22_y4, x23_y4, x24_y4, x25_y4, x26_y4, x27_y4, x28_y4, x29_y4, x30_y4, x31_y4, x32_y4, x33_y4, x34_y4, x35_y4, x36_y4, x37_y4, x38_y4, x39_y4, x40_y4, x41_y4, x42_y4, x43_y4, x44_y4, x45_y4, x46_y4, x47_y4, x48_y4, x49_y4, x50_y4, x51_y4, x52_y4, x53_y4, x54_y4, x55_y4, x56_y4, x57_y4, x58_y4, x59_y4, x60_y4, x61_y4, x0_y5, x1_y5, x2_y5, x3_y5, x4_y5, x5_y5, x6_y5, x7_y5, x8_y5, x9_y5, x10_y5, x11_y5, x12_y5, x13_y5, x14_y5, x15_y5, x16_y5, x17_y5, x18_y5, x19_y5, x20_y5, x21_y5, x22_y5, x23_y5, x24_y5, x25_y5, x26_y5, x27_y5, x28_y5, x29_y5, x30_y5, x31_y5, x32_y5, x33_y5, x34_y5, x35_y5, x36_y5, x37_y5, x38_y5, x39_y5, x40_y5, x41_y5, x42_y5, x43_y5, x44_y5, x45_y5, x46_y5, x47_y5, x48_y5, x49_y5, x50_y5, x51_y5, x52_y5, x53_y5, x54_y5, x55_y5, x56_y5, x57_y5, x58_y5, x59_y5, x60_y5, x61_y5, x0_y6, x1_y6, x2_y6, x3_y6, x4_y6, x5_y6, x6_y6, x7_y6, x8_y6, x9_y6, x10_y6, x11_y6, x12_y6, x13_y6, x14_y6, x15_y6, x16_y6, x17_y6, x18_y6, x19_y6, x20_y6, x21_y6, x22_y6, x23_y6, x24_y6, x25_y6, x26_y6, x27_y6, x28_y6, x29_y6, x30_y6, x31_y6, x32_y6, x33_y6, x34_y6, x35_y6, x36_y6, x37_y6, x38_y6, x39_y6, x40_y6, x41_y6, x42_y6, x43_y6, x44_y6, x45_y6, x46_y6, x47_y6, x48_y6, x49_y6, x50_y6, x51_y6, x52_y6, x53_y6, x54_y6, x55_y6, x56_y6, x57_y6, x58_y6, x59_y6, x60_y6, x61_y6, x0_y7, x1_y7, x2_y7, x3_y7, x4_y7, x5_y7, x6_y7, x7_y7, x8_y7, x9_y7, x10_y7, x11_y7, x12_y7, x13_y7, x14_y7, x15_y7, x16_y7, x17_y7, x18_y7, x19_y7, x20_y7, x21_y7, x22_y7, x23_y7, x24_y7, x25_y7, x26_y7, x27_y7, x28_y7, x29_y7, x30_y7, x31_y7, x32_y7, x33_y7, x34_y7, x35_y7, x36_y7, x37_y7, x38_y7, x39_y7, x40_y7, x41_y7, x42_y7, x43_y7, x44_y7, x45_y7, x46_y7, x47_y7, x48_y7, x49_y7, x50_y7, x51_y7, x52_y7, x53_y7, x54_y7, x55_y7, x56_y7, x57_y7, x58_y7, x59_y7, x60_y7, x61_y7, x0_y8, x1_y8, x2_y8, x3_y8, x4_y8, x5_y8, x6_y8, x7_y8, x8_y8, x9_y8, x10_y8, x11_y8, x12_y8, x13_y8, x14_y8, x15_y8, x16_y8, x17_y8, x18_y8, x19_y8, x20_y8, x21_y8, x22_y8, x23_y8, x24_y8, x25_y8, x26_y8, x27_y8, x28_y8, x29_y8, x30_y8, x31_y8, x32_y8, x33_y8, x34_y8, x35_y8, x36_y8, x37_y8, x38_y8, x39_y8, x40_y8, x41_y8, x42_y8, x43_y8, x44_y8, x45_y8, x46_y8, x47_y8, x48_y8, x49_y8, x50_y8, x51_y8, x52_y8, x53_y8, x54_y8, x55_y8, x56_y8, x57_y8, x58_y8, x59_y8, x60_y8, x61_y8, x0_y9, x1_y9, x2_y9, x3_y9, x4_y9, x5_y9, x6_y9, x7_y9, x8_y9, x9_y9, x10_y9, x11_y9, x12_y9, x13_y9, x14_y9, x15_y9, x16_y9, x17_y9, x18_y9, x19_y9, x20_y9, x21_y9, x22_y9, x23_y9, x24_y9, x25_y9, x26_y9, x27_y9, x28_y9, x29_y9, x30_y9, x31_y9, x32_y9, x33_y9, x34_y9, x35_y9, x36_y9, x37_y9, x38_y9, x39_y9, x40_y9, x41_y9, x42_y9, x43_y9, x44_y9, x45_y9, x46_y9, x47_y9, x48_y9, x49_y9, x50_y9, x51_y9, x52_y9, x53_y9, x54_y9, x55_y9, x56_y9, x57_y9, x58_y9, x59_y9, x60_y9, x61_y9, x0_y10, x1_y10, x2_y10, x3_y10, x4_y10, x5_y10, x6_y10, x7_y10, x8_y10, x9_y10, x10_y10, x11_y10, x12_y10, x13_y10, x14_y10, x15_y10, x16_y10, x17_y10, x18_y10, x19_y10, x20_y10, x21_y10, x22_y10, x23_y10, x24_y10, x25_y10, x26_y10, x27_y10, x28_y10, x29_y10, x30_y10, x31_y10, x32_y10, x33_y10, x34_y10, x35_y10, x36_y10, x37_y10, x38_y10, x39_y10, x40_y10, x41_y10, x42_y10, x43_y10, x44_y10, x45_y10, x46_y10, x47_y10, x48_y10, x49_y10, x50_y10, x51_y10, x52_y10, x53_y10, x54_y10, x55_y10, x56_y10, x57_y10, x58_y10, x59_y10, x60_y10, x61_y10, x0_y11, x1_y11, x2_y11, x3_y11, x4_y11, x5_y11, x6_y11, x7_y11, x8_y11, x9_y11, x10_y11, x11_y11, x12_y11, x13_y11, x14_y11, x15_y11, x16_y11, x17_y11, x18_y11, x19_y11, x20_y11, x21_y11, x22_y11, x23_y11, x24_y11, x25_y11, x26_y11, x27_y11, x28_y11, x29_y11, x30_y11, x31_y11, x32_y11, x33_y11, x34_y11, x35_y11, x36_y11, x37_y11, x38_y11, x39_y11, x40_y11, x41_y11, x42_y11, x43_y11, x44_y11, x45_y11, x46_y11, x47_y11, x48_y11, x49_y11, x50_y11, x51_y11, x52_y11, x53_y11, x54_y11, x55_y11, x56_y11, x57_y11, x58_y11, x59_y11, x60_y11, x61_y11, x0_y12, x1_y12, x2_y12, x3_y12, x4_y12, x5_y12, x6_y12, x7_y12, x8_y12, x9_y12, x10_y12, x11_y12, x12_y12, x13_y12, x14_y12, x15_y12, x16_y12, x17_y12, x18_y12, x19_y12, x20_y12, x21_y12, x22_y12, x23_y12, x24_y12, x25_y12, x26_y12, x27_y12, x28_y12, x29_y12, x30_y12, x31_y12, x32_y12, x33_y12, x34_y12, x35_y12, x36_y12, x37_y12, x38_y12, x39_y12, x40_y12, x41_y12, x42_y12, x43_y12, x44_y12, x45_y12, x46_y12, x47_y12, x48_y12, x49_y12, x50_y12, x51_y12, x52_y12, x53_y12, x54_y12, x55_y12, x56_y12, x57_y12, x58_y12, x59_y12, x60_y12, x61_y12, x0_y13, x1_y13, x2_y13, x3_y13, x4_y13, x5_y13, x6_y13, x7_y13, x8_y13, x9_y13, x10_y13, x11_y13, x12_y13, x13_y13, x14_y13, x15_y13, x16_y13, x17_y13, x18_y13, x19_y13, x20_y13, x21_y13, x22_y13, x23_y13, x24_y13, x25_y13, x26_y13, x27_y13, x28_y13, x29_y13, x30_y13, x31_y13, x32_y13, x33_y13, x34_y13, x35_y13, x36_y13, x37_y13, x38_y13, x39_y13, x40_y13, x41_y13, x42_y13, x43_y13, x44_y13, x45_y13, x46_y13, x47_y13, x48_y13, x49_y13, x50_y13, x51_y13, x52_y13, x53_y13, x54_y13, x55_y13, x56_y13, x57_y13, x58_y13, x59_y13, x60_y13, x61_y13, x0_y14, x1_y14, x2_y14, x3_y14, x4_y14, x5_y14, x6_y14, x7_y14, x8_y14, x9_y14, x10_y14, x11_y14, x12_y14, x13_y14, x14_y14, x15_y14, x16_y14, x17_y14, x18_y14, x19_y14, x20_y14, x21_y14, x22_y14, x23_y14, x24_y14, x25_y14, x26_y14, x27_y14, x28_y14, x29_y14, x30_y14, x31_y14, x32_y14, x33_y14, x34_y14, x35_y14, x36_y14, x37_y14, x38_y14, x39_y14, x40_y14, x41_y14, x42_y14, x43_y14, x44_y14, x45_y14, x46_y14, x47_y14, x48_y14, x49_y14, x50_y14, x51_y14, x52_y14, x53_y14, x54_y14, x55_y14, x56_y14, x57_y14, x58_y14, x59_y14, x60_y14, x61_y14, x0_y15, x1_y15, x2_y15, x3_y15, x4_y15, x5_y15, x6_y15, x7_y15, x8_y15, x9_y15, x10_y15, x11_y15, x12_y15, x13_y15, x14_y15, x15_y15, x16_y15, x17_y15, x18_y15, x19_y15, x20_y15, x21_y15, x22_y15, x23_y15, x24_y15, x25_y15, x26_y15, x27_y15, x28_y15, x29_y15, x30_y15, x31_y15, x32_y15, x33_y15, x34_y15, x35_y15, x36_y15, x37_y15, x38_y15, x39_y15, x40_y15, x41_y15, x42_y15, x43_y15, x44_y15, x45_y15, x46_y15, x47_y15, x48_y15, x49_y15, x50_y15, x51_y15, x52_y15, x53_y15, x54_y15, x55_y15, x56_y15, x57_y15, x58_y15, x59_y15, x60_y15, x61_y15, x0_y16, x1_y16, x2_y16, x3_y16, x4_y16, x5_y16, x6_y16, x7_y16, x8_y16, x9_y16, x10_y16, x11_y16, x12_y16, x13_y16, x14_y16, x15_y16, x16_y16, x17_y16, x18_y16, x19_y16, x20_y16, x21_y16, x22_y16, x23_y16, x24_y16, x25_y16, x26_y16, x27_y16, x28_y16, x29_y16, x30_y16, x31_y16, x32_y16, x33_y16, x34_y16, x35_y16, x36_y16, x37_y16, x38_y16, x39_y16, x40_y16, x41_y16, x42_y16, x43_y16, x44_y16, x45_y16, x46_y16, x47_y16, x48_y16, x49_y16, x50_y16, x51_y16, x52_y16, x53_y16, x54_y16, x55_y16, x56_y16, x57_y16, x58_y16, x59_y16, x60_y16, x61_y16, x0_y17, x1_y17, x2_y17, x3_y17, x4_y17, x5_y17, x6_y17, x7_y17, x8_y17, x9_y17, x10_y17, x11_y17, x12_y17, x13_y17, x14_y17, x15_y17, x16_y17, x17_y17, x18_y17, x19_y17, x20_y17, x21_y17, x22_y17, x23_y17, x24_y17, x25_y17, x26_y17, x27_y17, x28_y17, x29_y17, x30_y17, x31_y17, x32_y17, x33_y17, x34_y17, x35_y17, x36_y17, x37_y17, x38_y17, x39_y17, x40_y17, x41_y17, x42_y17, x43_y17, x44_y17, x45_y17, x46_y17, x47_y17, x48_y17, x49_y17, x50_y17, x51_y17, x52_y17, x53_y17, x54_y17, x55_y17, x56_y17, x57_y17, x58_y17, x59_y17, x60_y17, x61_y17, x0_y18, x1_y18, x2_y18, x3_y18, x4_y18, x5_y18, x6_y18, x7_y18, x8_y18, x9_y18, x10_y18, x11_y18, x12_y18, x13_y18, x14_y18, x15_y18, x16_y18, x17_y18, x18_y18, x19_y18, x20_y18, x21_y18, x22_y18, x23_y18, x24_y18, x25_y18, x26_y18, x27_y18, x28_y18, x29_y18, x30_y18, x31_y18, x32_y18, x33_y18, x34_y18, x35_y18, x36_y18, x37_y18, x38_y18, x39_y18, x40_y18, x41_y18, x42_y18, x43_y18, x44_y18, x45_y18, x46_y18, x47_y18, x48_y18, x49_y18, x50_y18, x51_y18, x52_y18, x53_y18, x54_y18, x55_y18, x56_y18, x57_y18, x58_y18, x59_y18, x60_y18, x61_y18, x0_y19, x1_y19, x2_y19, x3_y19, x4_y19, x5_y19, x6_y19, x7_y19, x8_y19, x9_y19, x10_y19, x11_y19, x12_y19, x13_y19, x14_y19, x15_y19, x16_y19, x17_y19, x18_y19, x19_y19, x20_y19, x21_y19, x22_y19, x23_y19, x24_y19, x25_y19, x26_y19, x27_y19, x28_y19, x29_y19, x30_y19, x31_y19, x32_y19, x33_y19, x34_y19, x35_y19, x36_y19, x37_y19, x38_y19, x39_y19, x40_y19, x41_y19, x42_y19, x43_y19, x44_y19, x45_y19, x46_y19, x47_y19, x48_y19, x49_y19, x50_y19, x51_y19, x52_y19, x53_y19, x54_y19, x55_y19, x56_y19, x57_y19, x58_y19, x59_y19, x60_y19, x61_y19, x0_y20, x1_y20, x2_y20, x3_y20, x4_y20, x5_y20, x6_y20, x7_y20, x8_y20, x9_y20, x10_y20, x11_y20, x12_y20, x13_y20, x14_y20, x15_y20, x16_y20, x17_y20, x18_y20, x19_y20, x20_y20, x21_y20, x22_y20, x23_y20, x24_y20, x25_y20, x26_y20, x27_y20, x28_y20, x29_y20, x30_y20, x31_y20, x32_y20, x33_y20, x34_y20, x35_y20, x36_y20, x37_y20, x38_y20, x39_y20, x40_y20, x41_y20, x42_y20, x43_y20, x44_y20, x45_y20, x46_y20, x47_y20, x48_y20, x49_y20, x50_y20, x51_y20, x52_y20, x53_y20, x54_y20, x55_y20, x56_y20, x57_y20, x58_y20, x59_y20, x60_y20, x61_y20, x0_y21, x1_y21, x2_y21, x3_y21, x4_y21, x5_y21, x6_y21, x7_y21, x8_y21, x9_y21, x10_y21, x11_y21, x12_y21, x13_y21, x14_y21, x15_y21, x16_y21, x17_y21, x18_y21, x19_y21, x20_y21, x21_y21, x22_y21, x23_y21, x24_y21, x25_y21, x26_y21, x27_y21, x28_y21, x29_y21, x30_y21, x31_y21, x32_y21, x33_y21, x34_y21, x35_y21, x36_y21, x37_y21, x38_y21, x39_y21, x40_y21, x41_y21, x42_y21, x43_y21, x44_y21, x45_y21, x46_y21, x47_y21, x48_y21, x49_y21, x50_y21, x51_y21, x52_y21, x53_y21, x54_y21, x55_y21, x56_y21, x57_y21, x58_y21, x59_y21, x60_y21, x61_y21, x0_y22, x1_y22, x2_y22, x3_y22, x4_y22, x5_y22, x6_y22, x7_y22, x8_y22, x9_y22, x10_y22, x11_y22, x12_y22, x13_y22, x14_y22, x15_y22, x16_y22, x17_y22, x18_y22, x19_y22, x20_y22, x21_y22, x22_y22, x23_y22, x24_y22, x25_y22, x26_y22, x27_y22, x28_y22, x29_y22, x30_y22, x31_y22, x32_y22, x33_y22, x34_y22, x35_y22, x36_y22, x37_y22, x38_y22, x39_y22, x40_y22, x41_y22, x42_y22, x43_y22, x44_y22, x45_y22, x46_y22, x47_y22, x48_y22, x49_y22, x50_y22, x51_y22, x52_y22, x53_y22, x54_y22, x55_y22, x56_y22, x57_y22, x58_y22, x59_y22, x60_y22, x61_y22, x0_y23, x1_y23, x2_y23, x3_y23, x4_y23, x5_y23, x6_y23, x7_y23, x8_y23, x9_y23, x10_y23, x11_y23, x12_y23, x13_y23, x14_y23, x15_y23, x16_y23, x17_y23, x18_y23, x19_y23, x20_y23, x21_y23, x22_y23, x23_y23, x24_y23, x25_y23, x26_y23, x27_y23, x28_y23, x29_y23, x30_y23, x31_y23, x32_y23, x33_y23, x34_y23, x35_y23, x36_y23, x37_y23, x38_y23, x39_y23, x40_y23, x41_y23, x42_y23, x43_y23, x44_y23, x45_y23, x46_y23, x47_y23, x48_y23, x49_y23, x50_y23, x51_y23, x52_y23, x53_y23, x54_y23, x55_y23, x56_y23, x57_y23, x58_y23, x59_y23, x60_y23, x61_y23, x0_y24, x1_y24, x2_y24, x3_y24, x4_y24, x5_y24, x6_y24, x7_y24, x8_y24, x9_y24, x10_y24, x11_y24, x12_y24, x13_y24, x14_y24, x15_y24, x16_y24, x17_y24, x18_y24, x19_y24, x20_y24, x21_y24, x22_y24, x23_y24, x24_y24, x25_y24, x26_y24, x27_y24, x28_y24, x29_y24, x30_y24, x31_y24, x32_y24, x33_y24, x34_y24, x35_y24, x36_y24, x37_y24, x38_y24, x39_y24, x40_y24, x41_y24, x42_y24, x43_y24, x44_y24, x45_y24, x46_y24, x47_y24, x48_y24, x49_y24, x50_y24, x51_y24, x52_y24, x53_y24, x54_y24, x55_y24, x56_y24, x57_y24, x58_y24, x59_y24, x60_y24, x61_y24, x0_y25, x1_y25, x2_y25, x3_y25, x4_y25, x5_y25, x6_y25, x7_y25, x8_y25, x9_y25, x10_y25, x11_y25, x12_y25, x13_y25, x14_y25, x15_y25, x16_y25, x17_y25, x18_y25, x19_y25, x20_y25, x21_y25, x22_y25, x23_y25, x24_y25, x25_y25, x26_y25, x27_y25, x28_y25, x29_y25, x30_y25, x31_y25, x32_y25, x33_y25, x34_y25, x35_y25, x36_y25, x37_y25, x38_y25, x39_y25, x40_y25, x41_y25, x42_y25, x43_y25, x44_y25, x45_y25, x46_y25, x47_y25, x48_y25, x49_y25, x50_y25, x51_y25, x52_y25, x53_y25, x54_y25, x55_y25, x56_y25, x57_y25, x58_y25, x59_y25, x60_y25, x61_y25, x0_y26, x1_y26, x2_y26, x3_y26, x4_y26, x5_y26, x6_y26, x7_y26, x8_y26, x9_y26, x10_y26, x11_y26, x12_y26, x13_y26, x14_y26, x15_y26, x16_y26, x17_y26, x18_y26, x19_y26, x20_y26, x21_y26, x22_y26, x23_y26, x24_y26, x25_y26, x26_y26, x27_y26, x28_y26, x29_y26, x30_y26, x31_y26, x32_y26, x33_y26, x34_y26, x35_y26, x36_y26, x37_y26, x38_y26, x39_y26, x40_y26, x41_y26, x42_y26, x43_y26, x44_y26, x45_y26, x46_y26, x47_y26, x48_y26, x49_y26, x50_y26, x51_y26, x52_y26, x53_y26, x54_y26, x55_y26, x56_y26, x57_y26, x58_y26, x59_y26, x60_y26, x61_y26, x0_y27, x1_y27, x2_y27, x3_y27, x4_y27, x5_y27, x6_y27, x7_y27, x8_y27, x9_y27, x10_y27, x11_y27, x12_y27, x13_y27, x14_y27, x15_y27, x16_y27, x17_y27, x18_y27, x19_y27, x20_y27, x21_y27, x22_y27, x23_y27, x24_y27, x25_y27, x26_y27, x27_y27, x28_y27, x29_y27, x30_y27, x31_y27, x32_y27, x33_y27, x34_y27, x35_y27, x36_y27, x37_y27, x38_y27, x39_y27, x40_y27, x41_y27, x42_y27, x43_y27, x44_y27, x45_y27, x46_y27, x47_y27, x48_y27, x49_y27, x50_y27, x51_y27, x52_y27, x53_y27, x54_y27, x55_y27, x56_y27, x57_y27, x58_y27, x59_y27, x60_y27, x61_y27, x0_y28, x1_y28, x2_y28, x3_y28, x4_y28, x5_y28, x6_y28, x7_y28, x8_y28, x9_y28, x10_y28, x11_y28, x12_y28, x13_y28, x14_y28, x15_y28, x16_y28, x17_y28, x18_y28, x19_y28, x20_y28, x21_y28, x22_y28, x23_y28, x24_y28, x25_y28, x26_y28, x27_y28, x28_y28, x29_y28, x30_y28, x31_y28, x32_y28, x33_y28, x34_y28, x35_y28, x36_y28, x37_y28, x38_y28, x39_y28, x40_y28, x41_y28, x42_y28, x43_y28, x44_y28, x45_y28, x46_y28, x47_y28, x48_y28, x49_y28, x50_y28, x51_y28, x52_y28, x53_y28, x54_y28, x55_y28, x56_y28, x57_y28, x58_y28, x59_y28, x60_y28, x61_y28, x0_y29, x1_y29, x2_y29, x3_y29, x4_y29, x5_y29, x6_y29, x7_y29, x8_y29, x9_y29, x10_y29, x11_y29, x12_y29, x13_y29, x14_y29, x15_y29, x16_y29, x17_y29, x18_y29, x19_y29, x20_y29, x21_y29, x22_y29, x23_y29, x24_y29, x25_y29, x26_y29, x27_y29, x28_y29, x29_y29, x30_y29, x31_y29, x32_y29, x33_y29, x34_y29, x35_y29, x36_y29, x37_y29, x38_y29, x39_y29, x40_y29, x41_y29, x42_y29, x43_y29, x44_y29, x45_y29, x46_y29, x47_y29, x48_y29, x49_y29, x50_y29, x51_y29, x52_y29, x53_y29, x54_y29, x55_y29, x56_y29, x57_y29, x58_y29, x59_y29, x60_y29, x61_y29, x0_y30, x1_y30, x2_y30, x3_y30, x4_y30, x5_y30, x6_y30, x7_y30, x8_y30, x9_y30, x10_y30, x11_y30, x12_y30, x13_y30, x14_y30, x15_y30, x16_y30, x17_y30, x18_y30, x19_y30, x20_y30, x21_y30, x22_y30, x23_y30, x24_y30, x25_y30, x26_y30, x27_y30, x28_y30, x29_y30, x30_y30, x31_y30, x32_y30, x33_y30, x34_y30, x35_y30, x36_y30, x37_y30, x38_y30, x39_y30, x40_y30, x41_y30, x42_y30, x43_y30, x44_y30, x45_y30, x46_y30, x47_y30, x48_y30, x49_y30, x50_y30, x51_y30, x52_y30, x53_y30, x54_y30, x55_y30, x56_y30, x57_y30, x58_y30, x59_y30, x60_y30, x61_y30, x0_y31, x1_y31, x2_y31, x3_y31, x4_y31, x5_y31, x6_y31, x7_y31, x8_y31, x9_y31, x10_y31, x11_y31, x12_y31, x13_y31, x14_y31, x15_y31, x16_y31, x17_y31, x18_y31, x19_y31, x20_y31, x21_y31, x22_y31, x23_y31, x24_y31, x25_y31, x26_y31, x27_y31, x28_y31, x29_y31, x30_y31, x31_y31, x32_y31, x33_y31, x34_y31, x35_y31, x36_y31, x37_y31, x38_y31, x39_y31, x40_y31, x41_y31, x42_y31, x43_y31, x44_y31, x45_y31, x46_y31, x47_y31, x48_y31, x49_y31, x50_y31, x51_y31, x52_y31, x53_y31, x54_y31, x55_y31, x56_y31, x57_y31, x58_y31, x59_y31, x60_y31, x61_y31, x0_y32, x1_y32, x2_y32, x3_y32, x4_y32, x5_y32, x6_y32, x7_y32, x8_y32, x9_y32, x10_y32, x11_y32, x12_y32, x13_y32, x14_y32, x15_y32, x16_y32, x17_y32, x18_y32, x19_y32, x20_y32, x21_y32, x22_y32, x23_y32, x24_y32, x25_y32, x26_y32, x27_y32, x28_y32, x29_y32, x30_y32, x31_y32, x32_y32, x33_y32, x34_y32, x35_y32, x36_y32, x37_y32, x38_y32, x39_y32, x40_y32, x41_y32, x42_y32, x43_y32, x44_y32, x45_y32, x46_y32, x47_y32, x48_y32, x49_y32, x50_y32, x51_y32, x52_y32, x53_y32, x54_y32, x55_y32, x56_y32, x57_y32, x58_y32, x59_y32, x60_y32, x61_y32, x0_y33, x1_y33, x2_y33, x3_y33, x4_y33, x5_y33, x6_y33, x7_y33, x8_y33, x9_y33, x10_y33, x11_y33, x12_y33, x13_y33, x14_y33, x15_y33, x16_y33, x17_y33, x18_y33, x19_y33, x20_y33, x21_y33, x22_y33, x23_y33, x24_y33, x25_y33, x26_y33, x27_y33, x28_y33, x29_y33, x30_y33, x31_y33, x32_y33, x33_y33, x34_y33, x35_y33, x36_y33, x37_y33, x38_y33, x39_y33, x40_y33, x41_y33, x42_y33, x43_y33, x44_y33, x45_y33, x46_y33, x47_y33, x48_y33, x49_y33, x50_y33, x51_y33, x52_y33, x53_y33, x54_y33, x55_y33, x56_y33, x57_y33, x58_y33, x59_y33, x60_y33, x61_y33, x0_y34, x1_y34, x2_y34, x3_y34, x4_y34, x5_y34, x6_y34, x7_y34, x8_y34, x9_y34, x10_y34, x11_y34, x12_y34, x13_y34, x14_y34, x15_y34, x16_y34, x17_y34, x18_y34, x19_y34, x20_y34, x21_y34, x22_y34, x23_y34, x24_y34, x25_y34, x26_y34, x27_y34, x28_y34, x29_y34, x30_y34, x31_y34, x32_y34, x33_y34, x34_y34, x35_y34, x36_y34, x37_y34, x38_y34, x39_y34, x40_y34, x41_y34, x42_y34, x43_y34, x44_y34, x45_y34, x46_y34, x47_y34, x48_y34, x49_y34, x50_y34, x51_y34, x52_y34, x53_y34, x54_y34, x55_y34, x56_y34, x57_y34, x58_y34, x59_y34, x60_y34, x61_y34, x0_y35, x1_y35, x2_y35, x3_y35, x4_y35, x5_y35, x6_y35, x7_y35, x8_y35, x9_y35, x10_y35, x11_y35, x12_y35, x13_y35, x14_y35, x15_y35, x16_y35, x17_y35, x18_y35, x19_y35, x20_y35, x21_y35, x22_y35, x23_y35, x24_y35, x25_y35, x26_y35, x27_y35, x28_y35, x29_y35, x30_y35, x31_y35, x32_y35, x33_y35, x34_y35, x35_y35, x36_y35, x37_y35, x38_y35, x39_y35, x40_y35, x41_y35, x42_y35, x43_y35, x44_y35, x45_y35, x46_y35, x47_y35, x48_y35, x49_y35, x50_y35, x51_y35, x52_y35, x53_y35, x54_y35, x55_y35, x56_y35, x57_y35, x58_y35, x59_y35, x60_y35, x61_y35, x0_y36, x1_y36, x2_y36, x3_y36, x4_y36, x5_y36, x6_y36, x7_y36, x8_y36, x9_y36, x10_y36, x11_y36, x12_y36, x13_y36, x14_y36, x15_y36, x16_y36, x17_y36, x18_y36, x19_y36, x20_y36, x21_y36, x22_y36, x23_y36, x24_y36, x25_y36, x26_y36, x27_y36, x28_y36, x29_y36, x30_y36, x31_y36, x32_y36, x33_y36, x34_y36, x35_y36, x36_y36, x37_y36, x38_y36, x39_y36, x40_y36, x41_y36, x42_y36, x43_y36, x44_y36, x45_y36, x46_y36, x47_y36, x48_y36, x49_y36, x50_y36, x51_y36, x52_y36, x53_y36, x54_y36, x55_y36, x56_y36, x57_y36, x58_y36, x59_y36, x60_y36, x61_y36, x0_y37, x1_y37, x2_y37, x3_y37, x4_y37, x5_y37, x6_y37, x7_y37, x8_y37, x9_y37, x10_y37, x11_y37, x12_y37, x13_y37, x14_y37, x15_y37, x16_y37, x17_y37, x18_y37, x19_y37, x20_y37, x21_y37, x22_y37, x23_y37, x24_y37, x25_y37, x26_y37, x27_y37, x28_y37, x29_y37, x30_y37, x31_y37, x32_y37, x33_y37, x34_y37, x35_y37, x36_y37, x37_y37, x38_y37, x39_y37, x40_y37, x41_y37, x42_y37, x43_y37, x44_y37, x45_y37, x46_y37, x47_y37, x48_y37, x49_y37, x50_y37, x51_y37, x52_y37, x53_y37, x54_y37, x55_y37, x56_y37, x57_y37, x58_y37, x59_y37, x60_y37, x61_y37, x0_y38, x1_y38, x2_y38, x3_y38, x4_y38, x5_y38, x6_y38, x7_y38, x8_y38, x9_y38, x10_y38, x11_y38, x12_y38, x13_y38, x14_y38, x15_y38, x16_y38, x17_y38, x18_y38, x19_y38, x20_y38, x21_y38, x22_y38, x23_y38, x24_y38, x25_y38, x26_y38, x27_y38, x28_y38, x29_y38, x30_y38, x31_y38, x32_y38, x33_y38, x34_y38, x35_y38, x36_y38, x37_y38, x38_y38, x39_y38, x40_y38, x41_y38, x42_y38, x43_y38, x44_y38, x45_y38, x46_y38, x47_y38, x48_y38, x49_y38, x50_y38, x51_y38, x52_y38, x53_y38, x54_y38, x55_y38, x56_y38, x57_y38, x58_y38, x59_y38, x60_y38, x61_y38, x0_y39, x1_y39, x2_y39, x3_y39, x4_y39, x5_y39, x6_y39, x7_y39, x8_y39, x9_y39, x10_y39, x11_y39, x12_y39, x13_y39, x14_y39, x15_y39, x16_y39, x17_y39, x18_y39, x19_y39, x20_y39, x21_y39, x22_y39, x23_y39, x24_y39, x25_y39, x26_y39, x27_y39, x28_y39, x29_y39, x30_y39, x31_y39, x32_y39, x33_y39, x34_y39, x35_y39, x36_y39, x37_y39, x38_y39, x39_y39, x40_y39, x41_y39, x42_y39, x43_y39, x44_y39, x45_y39, x46_y39, x47_y39, x48_y39, x49_y39, x50_y39, x51_y39, x52_y39, x53_y39, x54_y39, x55_y39, x56_y39, x57_y39, x58_y39, x59_y39, x60_y39, x61_y39, x0_y40, x1_y40, x2_y40, x3_y40, x4_y40, x5_y40, x6_y40, x7_y40, x8_y40, x9_y40, x10_y40, x11_y40, x12_y40, x13_y40, x14_y40, x15_y40, x16_y40, x17_y40, x18_y40, x19_y40, x20_y40, x21_y40, x22_y40, x23_y40, x24_y40, x25_y40, x26_y40, x27_y40, x28_y40, x29_y40, x30_y40, x31_y40, x32_y40, x33_y40, x34_y40, x35_y40, x36_y40, x37_y40, x38_y40, x39_y40, x40_y40, x41_y40, x42_y40, x43_y40, x44_y40, x45_y40, x46_y40, x47_y40, x48_y40, x49_y40, x50_y40, x51_y40, x52_y40, x53_y40, x54_y40, x55_y40, x56_y40, x57_y40, x58_y40, x59_y40, x60_y40, x61_y40, x0_y41, x1_y41, x2_y41, x3_y41, x4_y41, x5_y41, x6_y41, x7_y41, x8_y41, x9_y41, x10_y41, x11_y41, x12_y41, x13_y41, x14_y41, x15_y41, x16_y41, x17_y41, x18_y41, x19_y41, x20_y41, x21_y41, x22_y41, x23_y41, x24_y41, x25_y41, x26_y41, x27_y41, x28_y41, x29_y41, x30_y41, x31_y41, x32_y41, x33_y41, x34_y41, x35_y41, x36_y41, x37_y41, x38_y41, x39_y41, x40_y41, x41_y41, x42_y41, x43_y41, x44_y41, x45_y41, x46_y41, x47_y41, x48_y41, x49_y41, x50_y41, x51_y41, x52_y41, x53_y41, x54_y41, x55_y41, x56_y41, x57_y41, x58_y41, x59_y41, x60_y41, x61_y41, x0_y42, x1_y42, x2_y42, x3_y42, x4_y42, x5_y42, x6_y42, x7_y42, x8_y42, x9_y42, x10_y42, x11_y42, x12_y42, x13_y42, x14_y42, x15_y42, x16_y42, x17_y42, x18_y42, x19_y42, x20_y42, x21_y42, x22_y42, x23_y42, x24_y42, x25_y42, x26_y42, x27_y42, x28_y42, x29_y42, x30_y42, x31_y42, x32_y42, x33_y42, x34_y42, x35_y42, x36_y42, x37_y42, x38_y42, x39_y42, x40_y42, x41_y42, x42_y42, x43_y42, x44_y42, x45_y42, x46_y42, x47_y42, x48_y42, x49_y42, x50_y42, x51_y42, x52_y42, x53_y42, x54_y42, x55_y42, x56_y42, x57_y42, x58_y42, x59_y42, x60_y42, x61_y42, x0_y43, x1_y43, x2_y43, x3_y43, x4_y43, x5_y43, x6_y43, x7_y43, x8_y43, x9_y43, x10_y43, x11_y43, x12_y43, x13_y43, x14_y43, x15_y43, x16_y43, x17_y43, x18_y43, x19_y43, x20_y43, x21_y43, x22_y43, x23_y43, x24_y43, x25_y43, x26_y43, x27_y43, x28_y43, x29_y43, x30_y43, x31_y43, x32_y43, x33_y43, x34_y43, x35_y43, x36_y43, x37_y43, x38_y43, x39_y43, x40_y43, x41_y43, x42_y43, x43_y43, x44_y43, x45_y43, x46_y43, x47_y43, x48_y43, x49_y43, x50_y43, x51_y43, x52_y43, x53_y43, x54_y43, x55_y43, x56_y43, x57_y43, x58_y43, x59_y43, x60_y43, x61_y43, x0_y44, x1_y44, x2_y44, x3_y44, x4_y44, x5_y44, x6_y44, x7_y44, x8_y44, x9_y44, x10_y44, x11_y44, x12_y44, x13_y44, x14_y44, x15_y44, x16_y44, x17_y44, x18_y44, x19_y44, x20_y44, x21_y44, x22_y44, x23_y44, x24_y44, x25_y44, x26_y44, x27_y44, x28_y44, x29_y44, x30_y44, x31_y44, x32_y44, x33_y44, x34_y44, x35_y44, x36_y44, x37_y44, x38_y44, x39_y44, x40_y44, x41_y44, x42_y44, x43_y44, x44_y44, x45_y44, x46_y44, x47_y44, x48_y44, x49_y44, x50_y44, x51_y44, x52_y44, x53_y44, x54_y44, x55_y44, x56_y44, x57_y44, x58_y44, x59_y44, x60_y44, x61_y44, x0_y45, x1_y45, x2_y45, x3_y45, x4_y45, x5_y45, x6_y45, x7_y45, x8_y45, x9_y45, x10_y45, x11_y45, x12_y45, x13_y45, x14_y45, x15_y45, x16_y45, x17_y45, x18_y45, x19_y45, x20_y45, x21_y45, x22_y45, x23_y45, x24_y45, x25_y45, x26_y45, x27_y45, x28_y45, x29_y45, x30_y45, x31_y45, x32_y45, x33_y45, x34_y45, x35_y45, x36_y45, x37_y45, x38_y45, x39_y45, x40_y45, x41_y45, x42_y45, x43_y45, x44_y45, x45_y45, x46_y45, x47_y45, x48_y45, x49_y45, x50_y45, x51_y45, x52_y45, x53_y45, x54_y45, x55_y45, x56_y45, x57_y45, x58_y45, x59_y45, x60_y45, x61_y45, x0_y46, x1_y46, x2_y46, x3_y46, x4_y46, x5_y46, x6_y46, x7_y46, x8_y46, x9_y46, x10_y46, x11_y46, x12_y46, x13_y46, x14_y46, x15_y46, x16_y46, x17_y46, x18_y46, x19_y46, x20_y46, x21_y46, x22_y46, x23_y46, x24_y46, x25_y46, x26_y46, x27_y46, x28_y46, x29_y46, x30_y46, x31_y46, x32_y46, x33_y46, x34_y46, x35_y46, x36_y46, x37_y46, x38_y46, x39_y46, x40_y46, x41_y46, x42_y46, x43_y46, x44_y46, x45_y46, x46_y46, x47_y46, x48_y46, x49_y46, x50_y46, x51_y46, x52_y46, x53_y46, x54_y46, x55_y46, x56_y46, x57_y46, x58_y46, x59_y46, x60_y46, x61_y46, x0_y47, x1_y47, x2_y47, x3_y47, x4_y47, x5_y47, x6_y47, x7_y47, x8_y47, x9_y47, x10_y47, x11_y47, x12_y47, x13_y47, x14_y47, x15_y47, x16_y47, x17_y47, x18_y47, x19_y47, x20_y47, x21_y47, x22_y47, x23_y47, x24_y47, x25_y47, x26_y47, x27_y47, x28_y47, x29_y47, x30_y47, x31_y47, x32_y47, x33_y47, x34_y47, x35_y47, x36_y47, x37_y47, x38_y47, x39_y47, x40_y47, x41_y47, x42_y47, x43_y47, x44_y47, x45_y47, x46_y47, x47_y47, x48_y47, x49_y47, x50_y47, x51_y47, x52_y47, x53_y47, x54_y47, x55_y47, x56_y47, x57_y47, x58_y47, x59_y47, x60_y47, x61_y47, x0_y48, x1_y48, x2_y48, x3_y48, x4_y48, x5_y48, x6_y48, x7_y48, x8_y48, x9_y48, x10_y48, x11_y48, x12_y48, x13_y48, x14_y48, x15_y48, x16_y48, x17_y48, x18_y48, x19_y48, x20_y48, x21_y48, x22_y48, x23_y48, x24_y48, x25_y48, x26_y48, x27_y48, x28_y48, x29_y48, x30_y48, x31_y48, x32_y48, x33_y48, x34_y48, x35_y48, x36_y48, x37_y48, x38_y48, x39_y48, x40_y48, x41_y48, x42_y48, x43_y48, x44_y48, x45_y48, x46_y48, x47_y48, x48_y48, x49_y48, x50_y48, x51_y48, x52_y48, x53_y48, x54_y48, x55_y48, x56_y48, x57_y48, x58_y48, x59_y48, x60_y48, x61_y48, x0_y49, x1_y49, x2_y49, x3_y49, x4_y49, x5_y49, x6_y49, x7_y49, x8_y49, x9_y49, x10_y49, x11_y49, x12_y49, x13_y49, x14_y49, x15_y49, x16_y49, x17_y49, x18_y49, x19_y49, x20_y49, x21_y49, x22_y49, x23_y49, x24_y49, x25_y49, x26_y49, x27_y49, x28_y49, x29_y49, x30_y49, x31_y49, x32_y49, x33_y49, x34_y49, x35_y49, x36_y49, x37_y49, x38_y49, x39_y49, x40_y49, x41_y49, x42_y49, x43_y49, x44_y49, x45_y49, x46_y49, x47_y49, x48_y49, x49_y49, x50_y49, x51_y49, x52_y49, x53_y49, x54_y49, x55_y49, x56_y49, x57_y49, x58_y49, x59_y49, x60_y49, x61_y49, x0_y50, x1_y50, x2_y50, x3_y50, x4_y50, x5_y50, x6_y50, x7_y50, x8_y50, x9_y50, x10_y50, x11_y50, x12_y50, x13_y50, x14_y50, x15_y50, x16_y50, x17_y50, x18_y50, x19_y50, x20_y50, x21_y50, x22_y50, x23_y50, x24_y50, x25_y50, x26_y50, x27_y50, x28_y50, x29_y50, x30_y50, x31_y50, x32_y50, x33_y50, x34_y50, x35_y50, x36_y50, x37_y50, x38_y50, x39_y50, x40_y50, x41_y50, x42_y50, x43_y50, x44_y50, x45_y50, x46_y50, x47_y50, x48_y50, x49_y50, x50_y50, x51_y50, x52_y50, x53_y50, x54_y50, x55_y50, x56_y50, x57_y50, x58_y50, x59_y50, x60_y50, x61_y50, x0_y51, x1_y51, x2_y51, x3_y51, x4_y51, x5_y51, x6_y51, x7_y51, x8_y51, x9_y51, x10_y51, x11_y51, x12_y51, x13_y51, x14_y51, x15_y51, x16_y51, x17_y51, x18_y51, x19_y51, x20_y51, x21_y51, x22_y51, x23_y51, x24_y51, x25_y51, x26_y51, x27_y51, x28_y51, x29_y51, x30_y51, x31_y51, x32_y51, x33_y51, x34_y51, x35_y51, x36_y51, x37_y51, x38_y51, x39_y51, x40_y51, x41_y51, x42_y51, x43_y51, x44_y51, x45_y51, x46_y51, x47_y51, x48_y51, x49_y51, x50_y51, x51_y51, x52_y51, x53_y51, x54_y51, x55_y51, x56_y51, x57_y51, x58_y51, x59_y51, x60_y51, x61_y51, x0_y52, x1_y52, x2_y52, x3_y52, x4_y52, x5_y52, x6_y52, x7_y52, x8_y52, x9_y52, x10_y52, x11_y52, x12_y52, x13_y52, x14_y52, x15_y52, x16_y52, x17_y52, x18_y52, x19_y52, x20_y52, x21_y52, x22_y52, x23_y52, x24_y52, x25_y52, x26_y52, x27_y52, x28_y52, x29_y52, x30_y52, x31_y52, x32_y52, x33_y52, x34_y52, x35_y52, x36_y52, x37_y52, x38_y52, x39_y52, x40_y52, x41_y52, x42_y52, x43_y52, x44_y52, x45_y52, x46_y52, x47_y52, x48_y52, x49_y52, x50_y52, x51_y52, x52_y52, x53_y52, x54_y52, x55_y52, x56_y52, x57_y52, x58_y52, x59_y52, x60_y52, x61_y52, x0_y53, x1_y53, x2_y53, x3_y53, x4_y53, x5_y53, x6_y53, x7_y53, x8_y53, x9_y53, x10_y53, x11_y53, x12_y53, x13_y53, x14_y53, x15_y53, x16_y53, x17_y53, x18_y53, x19_y53, x20_y53, x21_y53, x22_y53, x23_y53, x24_y53, x25_y53, x26_y53, x27_y53, x28_y53, x29_y53, x30_y53, x31_y53, x32_y53, x33_y53, x34_y53, x35_y53, x36_y53, x37_y53, x38_y53, x39_y53, x40_y53, x41_y53, x42_y53, x43_y53, x44_y53, x45_y53, x46_y53, x47_y53, x48_y53, x49_y53, x50_y53, x51_y53, x52_y53, x53_y53, x54_y53, x55_y53, x56_y53, x57_y53, x58_y53, x59_y53, x60_y53, x61_y53, x0_y54, x1_y54, x2_y54, x3_y54, x4_y54, x5_y54, x6_y54, x7_y54, x8_y54, x9_y54, x10_y54, x11_y54, x12_y54, x13_y54, x14_y54, x15_y54, x16_y54, x17_y54, x18_y54, x19_y54, x20_y54, x21_y54, x22_y54, x23_y54, x24_y54, x25_y54, x26_y54, x27_y54, x28_y54, x29_y54, x30_y54, x31_y54, x32_y54, x33_y54, x34_y54, x35_y54, x36_y54, x37_y54, x38_y54, x39_y54, x40_y54, x41_y54, x42_y54, x43_y54, x44_y54, x45_y54, x46_y54, x47_y54, x48_y54, x49_y54, x50_y54, x51_y54, x52_y54, x53_y54, x54_y54, x55_y54, x56_y54, x57_y54, x58_y54, x59_y54, x60_y54, x61_y54, x0_y55, x1_y55, x2_y55, x3_y55, x4_y55, x5_y55, x6_y55, x7_y55, x8_y55, x9_y55, x10_y55, x11_y55, x12_y55, x13_y55, x14_y55, x15_y55, x16_y55, x17_y55, x18_y55, x19_y55, x20_y55, x21_y55, x22_y55, x23_y55, x24_y55, x25_y55, x26_y55, x27_y55, x28_y55, x29_y55, x30_y55, x31_y55, x32_y55, x33_y55, x34_y55, x35_y55, x36_y55, x37_y55, x38_y55, x39_y55, x40_y55, x41_y55, x42_y55, x43_y55, x44_y55, x45_y55, x46_y55, x47_y55, x48_y55, x49_y55, x50_y55, x51_y55, x52_y55, x53_y55, x54_y55, x55_y55, x56_y55, x57_y55, x58_y55, x59_y55, x60_y55, x61_y55, x0_y56, x1_y56, x2_y56, x3_y56, x4_y56, x5_y56, x6_y56, x7_y56, x8_y56, x9_y56, x10_y56, x11_y56, x12_y56, x13_y56, x14_y56, x15_y56, x16_y56, x17_y56, x18_y56, x19_y56, x20_y56, x21_y56, x22_y56, x23_y56, x24_y56, x25_y56, x26_y56, x27_y56, x28_y56, x29_y56, x30_y56, x31_y56, x32_y56, x33_y56, x34_y56, x35_y56, x36_y56, x37_y56, x38_y56, x39_y56, x40_y56, x41_y56, x42_y56, x43_y56, x44_y56, x45_y56, x46_y56, x47_y56, x48_y56, x49_y56, x50_y56, x51_y56, x52_y56, x53_y56, x54_y56, x55_y56, x56_y56, x57_y56, x58_y56, x59_y56, x60_y56, x61_y56, x0_y57, x1_y57, x2_y57, x3_y57, x4_y57, x5_y57, x6_y57, x7_y57, x8_y57, x9_y57, x10_y57, x11_y57, x12_y57, x13_y57, x14_y57, x15_y57, x16_y57, x17_y57, x18_y57, x19_y57, x20_y57, x21_y57, x22_y57, x23_y57, x24_y57, x25_y57, x26_y57, x27_y57, x28_y57, x29_y57, x30_y57, x31_y57, x32_y57, x33_y57, x34_y57, x35_y57, x36_y57, x37_y57, x38_y57, x39_y57, x40_y57, x41_y57, x42_y57, x43_y57, x44_y57, x45_y57, x46_y57, x47_y57, x48_y57, x49_y57, x50_y57, x51_y57, x52_y57, x53_y57, x54_y57, x55_y57, x56_y57, x57_y57, x58_y57, x59_y57, x60_y57, x61_y57, x0_y58, x1_y58, x2_y58, x3_y58, x4_y58, x5_y58, x6_y58, x7_y58, x8_y58, x9_y58, x10_y58, x11_y58, x12_y58, x13_y58, x14_y58, x15_y58, x16_y58, x17_y58, x18_y58, x19_y58, x20_y58, x21_y58, x22_y58, x23_y58, x24_y58, x25_y58, x26_y58, x27_y58, x28_y58, x29_y58, x30_y58, x31_y58, x32_y58, x33_y58, x34_y58, x35_y58, x36_y58, x37_y58, x38_y58, x39_y58, x40_y58, x41_y58, x42_y58, x43_y58, x44_y58, x45_y58, x46_y58, x47_y58, x48_y58, x49_y58, x50_y58, x51_y58, x52_y58, x53_y58, x54_y58, x55_y58, x56_y58, x57_y58, x58_y58, x59_y58, x60_y58, x61_y58, x0_y59, x1_y59, x2_y59, x3_y59, x4_y59, x5_y59, x6_y59, x7_y59, x8_y59, x9_y59, x10_y59, x11_y59, x12_y59, x13_y59, x14_y59, x15_y59, x16_y59, x17_y59, x18_y59, x19_y59, x20_y59, x21_y59, x22_y59, x23_y59, x24_y59, x25_y59, x26_y59, x27_y59, x28_y59, x29_y59, x30_y59, x31_y59, x32_y59, x33_y59, x34_y59, x35_y59, x36_y59, x37_y59, x38_y59, x39_y59, x40_y59, x41_y59, x42_y59, x43_y59, x44_y59, x45_y59, x46_y59, x47_y59, x48_y59, x49_y59, x50_y59, x51_y59, x52_y59, x53_y59, x54_y59, x55_y59, x56_y59, x57_y59, x58_y59, x59_y59, x60_y59, x61_y59, x0_y60, x1_y60, x2_y60, x3_y60, x4_y60, x5_y60, x6_y60, x7_y60, x8_y60, x9_y60, x10_y60, x11_y60, x12_y60, x13_y60, x14_y60, x15_y60, x16_y60, x17_y60, x18_y60, x19_y60, x20_y60, x21_y60, x22_y60, x23_y60, x24_y60, x25_y60, x26_y60, x27_y60, x28_y60, x29_y60, x30_y60, x31_y60, x32_y60, x33_y60, x34_y60, x35_y60, x36_y60, x37_y60, x38_y60, x39_y60, x40_y60, x41_y60, x42_y60, x43_y60, x44_y60, x45_y60, x46_y60, x47_y60, x48_y60, x49_y60, x50_y60, x51_y60, x52_y60, x53_y60, x54_y60, x55_y60, x56_y60, x57_y60, x58_y60, x59_y60, x60_y60, x61_y60, x0_y61, x1_y61, x2_y61, x3_y61, x4_y61, x5_y61, x6_y61, x7_y61, x8_y61, x9_y61, x10_y61, x11_y61, x12_y61, x13_y61, x14_y61, x15_y61, x16_y61, x17_y61, x18_y61, x19_y61, x20_y61, x21_y61, x22_y61, x23_y61, x24_y61, x25_y61, x26_y61, x27_y61, x28_y61, x29_y61, x30_y61, x31_y61, x32_y61, x33_y61, x34_y61, x35_y61, x36_y61, x37_y61, x38_y61, x39_y61, x40_y61, x41_y61, x42_y61, x43_y61, x44_y61, x45_y61, x46_y61, x47_y61, x48_y61, x49_y61, x50_y61, x51_y61, x52_y61, x53_y61, x54_y61, x55_y61, x56_y61, x57_y61, x58_y61, x59_y61, x60_y61, x61_y61, x0_y62, x1_y62, x2_y62, x3_y62, x4_y62, x5_y62, x6_y62, x7_y62, x8_y62, x9_y62, x10_y62, x11_y62, x12_y62, x13_y62, x14_y62, x15_y62, x16_y62, x17_y62, x18_y62, x19_y62, x20_y62, x21_y62, x22_y62, x23_y62, x24_y62, x25_y62, x26_y62, x27_y62, x28_y62, x29_y62, x30_y62, x31_y62, x32_y62, x33_y62, x34_y62, x35_y62, x36_y62, x37_y62, x38_y62, x39_y62, x40_y62, x41_y62, x42_y62, x43_y62, x44_y62, x45_y62, x46_y62, x47_y62, x48_y62, x49_y62, x50_y62, x51_y62, x52_y62, x53_y62, x54_y62, x55_y62, x56_y62, x57_y62, x58_y62, x59_y62, x60_y62, x61_y62, x0_y63, x1_y63, x2_y63, x3_y63, x4_y63, x5_y63, x6_y63, x7_y63, x8_y63, x9_y63, x10_y63, x11_y63, x12_y63, x13_y63, x14_y63, x15_y63, x16_y63, x17_y63, x18_y63, x19_y63, x20_y63, x21_y63, x22_y63, x23_y63, x24_y63, x25_y63, x26_y63, x27_y63, x28_y63, x29_y63, x30_y63;


(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100100110001)
) lut_0_0 (
    .O(x0_y0),
    .I0(in4),
    .I1(in0),
    .I2(1'b0),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010110101011)
) lut_1_0 (
    .O(x1_y0),
    .I0(in0),
    .I1(1'b0),
    .I2(in4),
    .I3(in3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011000110111)
) lut_2_0 (
    .O(x2_y0),
    .I0(1'b0),
    .I1(1'b0),
    .I2(in2),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010101000011)
) lut_3_0 (
    .O(x3_y0),
    .I0(1'b0),
    .I1(1'b0),
    .I2(in0),
    .I3(x1_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111001101001)
) lut_4_0 (
    .O(x4_y0),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x1_y1),
    .I3(x2_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011001101010)
) lut_5_0 (
    .O(x5_y0),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x2_y2),
    .I3(x2_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010000010110)
) lut_6_0 (
    .O(x6_y0),
    .I0(1'b0),
    .I1(x3_y0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011010111000)
) lut_7_0 (
    .O(x7_y0),
    .I0(x5_y0),
    .I1(x5_y0),
    .I2(x5_y2),
    .I3(x5_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100010100111)
) lut_8_0 (
    .O(x8_y0),
    .I0(x5_y1),
    .I1(x6_y0),
    .I2(x6_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110101111100)
) lut_9_0 (
    .O(x9_y0),
    .I0(x7_y0),
    .I1(x6_y0),
    .I2(x6_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101110110010)
) lut_10_0 (
    .O(x10_y0),
    .I0(x8_y5),
    .I1(x7_y4),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111110111010)
) lut_11_0 (
    .O(x11_y0),
    .I0(x9_y0),
    .I1(x9_y0),
    .I2(1'b0),
    .I3(x9_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011010010010)
) lut_12_0 (
    .O(x12_y0),
    .I0(1'b0),
    .I1(x10_y5),
    .I2(1'b0),
    .I3(x10_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011000010011)
) lut_13_0 (
    .O(x13_y0),
    .I0(x11_y2),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101100101101)
) lut_14_0 (
    .O(x14_y0),
    .I0(x11_y0),
    .I1(x11_y0),
    .I2(x11_y0),
    .I3(x12_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110101110110)
) lut_15_0 (
    .O(x15_y0),
    .I0(x13_y0),
    .I1(1'b0),
    .I2(x13_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100111001000)
) lut_16_0 (
    .O(x16_y0),
    .I0(x13_y5),
    .I1(1'b0),
    .I2(x13_y0),
    .I3(x13_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011011111001)
) lut_17_0 (
    .O(x17_y0),
    .I0(x14_y1),
    .I1(x15_y0),
    .I2(x15_y0),
    .I3(x15_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001010010101)
) lut_18_0 (
    .O(x18_y0),
    .I0(x15_y0),
    .I1(x15_y5),
    .I2(x16_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111011110010)
) lut_19_0 (
    .O(x19_y0),
    .I0(x16_y4),
    .I1(1'b0),
    .I2(x17_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111011001001)
) lut_20_0 (
    .O(x20_y0),
    .I0(x17_y1),
    .I1(x17_y0),
    .I2(x18_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010110110111)
) lut_21_0 (
    .O(x21_y0),
    .I0(1'b0),
    .I1(x18_y0),
    .I2(1'b0),
    .I3(x19_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100001001011)
) lut_22_0 (
    .O(x22_y0),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x20_y0),
    .I3(x20_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110101101010)
) lut_23_0 (
    .O(x23_y0),
    .I0(1'b0),
    .I1(x21_y4),
    .I2(x20_y0),
    .I3(x20_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101001010111)
) lut_24_0 (
    .O(x24_y0),
    .I0(1'b0),
    .I1(x21_y0),
    .I2(x21_y0),
    .I3(x22_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111100110111)
) lut_25_0 (
    .O(x25_y0),
    .I0(x23_y5),
    .I1(x23_y2),
    .I2(x22_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111111000001)
) lut_26_0 (
    .O(x26_y0),
    .I0(x23_y0),
    .I1(x24_y0),
    .I2(1'b0),
    .I3(x24_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001011110111)
) lut_27_0 (
    .O(x27_y0),
    .I0(x25_y0),
    .I1(1'b0),
    .I2(x24_y2),
    .I3(x24_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110000100010)
) lut_28_0 (
    .O(x28_y0),
    .I0(1'b0),
    .I1(x26_y0),
    .I2(x26_y0),
    .I3(x25_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100111100101)
) lut_29_0 (
    .O(x29_y0),
    .I0(1'b0),
    .I1(x26_y0),
    .I2(x26_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101110000101)
) lut_30_0 (
    .O(x30_y0),
    .I0(1'b0),
    .I1(x28_y3),
    .I2(1'b0),
    .I3(x27_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001011111101)
) lut_31_0 (
    .O(x31_y0),
    .I0(x28_y0),
    .I1(x29_y1),
    .I2(x28_y0),
    .I3(x28_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010011010011)
) lut_32_0 (
    .O(x32_y0),
    .I0(x29_y0),
    .I1(x30_y1),
    .I2(x30_y5),
    .I3(x30_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011011100101)
) lut_33_0 (
    .O(x33_y0),
    .I0(x31_y2),
    .I1(1'b0),
    .I2(x31_y0),
    .I3(x30_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110110101100)
) lut_34_0 (
    .O(x34_y0),
    .I0(x32_y3),
    .I1(1'b0),
    .I2(x31_y1),
    .I3(x31_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010100111110)
) lut_35_0 (
    .O(x35_y0),
    .I0(x33_y2),
    .I1(x33_y0),
    .I2(x33_y0),
    .I3(x33_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001011000110)
) lut_36_0 (
    .O(x36_y0),
    .I0(x33_y3),
    .I1(x34_y0),
    .I2(x34_y3),
    .I3(x34_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001111001001)
) lut_37_0 (
    .O(x37_y0),
    .I0(x34_y0),
    .I1(x34_y0),
    .I2(x34_y3),
    .I3(x34_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110010100001)
) lut_38_0 (
    .O(x38_y0),
    .I0(x35_y0),
    .I1(x36_y0),
    .I2(x36_y0),
    .I3(x36_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000110100011)
) lut_39_0 (
    .O(x39_y0),
    .I0(x36_y4),
    .I1(x37_y2),
    .I2(x36_y0),
    .I3(x36_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001100101011)
) lut_40_0 (
    .O(x40_y0),
    .I0(x37_y0),
    .I1(x38_y4),
    .I2(1'b0),
    .I3(x37_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011100011110)
) lut_41_0 (
    .O(x41_y0),
    .I0(1'b0),
    .I1(x39_y2),
    .I2(x39_y0),
    .I3(x39_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100101001000)
) lut_42_0 (
    .O(x42_y0),
    .I0(1'b0),
    .I1(x39_y1),
    .I2(x39_y2),
    .I3(x40_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110010110101)
) lut_43_0 (
    .O(x43_y0),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x41_y0),
    .I3(x41_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010111010001)
) lut_44_0 (
    .O(x44_y0),
    .I0(x41_y0),
    .I1(1'b0),
    .I2(x41_y2),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010110101011)
) lut_45_0 (
    .O(x45_y0),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x43_y2),
    .I3(x43_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110010101110)
) lut_46_0 (
    .O(x46_y0),
    .I0(x44_y4),
    .I1(1'b0),
    .I2(x43_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011011001101)
) lut_47_0 (
    .O(x47_y0),
    .I0(x44_y0),
    .I1(1'b0),
    .I2(x44_y0),
    .I3(x44_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110111000001)
) lut_48_0 (
    .O(x48_y0),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x46_y2),
    .I3(x45_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111001010111)
) lut_49_0 (
    .O(x49_y0),
    .I0(1'b0),
    .I1(x47_y0),
    .I2(x47_y4),
    .I3(x46_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010000011000)
) lut_50_0 (
    .O(x50_y0),
    .I0(x47_y0),
    .I1(x47_y5),
    .I2(1'b0),
    .I3(x47_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011000100000)
) lut_51_0 (
    .O(x51_y0),
    .I0(1'b0),
    .I1(x49_y2),
    .I2(1'b0),
    .I3(x48_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100011100100)
) lut_52_0 (
    .O(x52_y0),
    .I0(x49_y0),
    .I1(x49_y0),
    .I2(x50_y1),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000000000001)
) lut_53_0 (
    .O(x53_y0),
    .I0(x50_y0),
    .I1(x50_y0),
    .I2(x50_y4),
    .I3(x50_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000101010101)
) lut_54_0 (
    .O(x54_y0),
    .I0(x52_y3),
    .I1(x51_y0),
    .I2(x52_y0),
    .I3(x51_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100111000000)
) lut_55_0 (
    .O(x55_y0),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x53_y2),
    .I3(x52_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110111011110)
) lut_56_0 (
    .O(x56_y0),
    .I0(1'b0),
    .I1(x54_y0),
    .I2(x53_y0),
    .I3(x54_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100010100010)
) lut_57_0 (
    .O(x57_y0),
    .I0(x54_y5),
    .I1(x54_y0),
    .I2(x55_y1),
    .I3(x55_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111010011111)
) lut_58_0 (
    .O(x58_y0),
    .I0(x55_y0),
    .I1(x56_y3),
    .I2(x56_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011010111110)
) lut_59_0 (
    .O(x59_y0),
    .I0(x57_y0),
    .I1(x56_y0),
    .I2(x56_y0),
    .I3(x57_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000000100011)
) lut_60_0 (
    .O(x60_y0),
    .I0(x57_y0),
    .I1(x58_y0),
    .I2(x57_y3),
    .I3(x57_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101111100000)
) lut_61_0 (
    .O(x61_y0),
    .I0(x59_y1),
    .I1(x59_y0),
    .I2(x59_y0),
    .I3(x59_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111110100001)
) lut_62_0 (
    .O(x62_y0),
    .I0(x60_y3),
    .I1(x59_y0),
    .I2(x59_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001101100101)
) lut_0_1 (
    .O(x0_y1),
    .I0(in0),
    .I1(1'b0),
    .I2(in0),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101100111011)
) lut_1_1 (
    .O(x1_y1),
    .I0(1'b0),
    .I1(in0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101001010111)
) lut_2_1 (
    .O(x2_y1),
    .I0(in0),
    .I1(in0),
    .I2(in4),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111010111110)
) lut_3_1 (
    .O(x3_y1),
    .I0(in0),
    .I1(in0),
    .I2(1'b0),
    .I3(x1_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100111101100)
) lut_4_1 (
    .O(x4_y1),
    .I0(x1_y2),
    .I1(x2_y0),
    .I2(x2_y5),
    .I3(x2_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101000010000)
) lut_5_1 (
    .O(x5_y1),
    .I0(1'b0),
    .I1(x2_y0),
    .I2(1'b0),
    .I3(x3_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100010111110)
) lut_6_1 (
    .O(x6_y1),
    .I0(x4_y3),
    .I1(x3_y0),
    .I2(x4_y0),
    .I3(x3_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111110110110)
) lut_7_1 (
    .O(x7_y1),
    .I0(x5_y0),
    .I1(x5_y0),
    .I2(1'b0),
    .I3(x4_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010000100110)
) lut_8_1 (
    .O(x8_y1),
    .I0(x6_y0),
    .I1(x5_y6),
    .I2(x6_y1),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001100110011)
) lut_9_1 (
    .O(x9_y1),
    .I0(x7_y5),
    .I1(x6_y6),
    .I2(x6_y1),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010100001001)
) lut_10_1 (
    .O(x10_y1),
    .I0(x8_y0),
    .I1(x7_y0),
    .I2(x7_y4),
    .I3(x8_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001001011110)
) lut_11_1 (
    .O(x11_y1),
    .I0(1'b0),
    .I1(x8_y3),
    .I2(1'b0),
    .I3(x9_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110101111111)
) lut_12_1 (
    .O(x12_y1),
    .I0(x10_y2),
    .I1(x9_y0),
    .I2(1'b0),
    .I3(x10_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000101111000)
) lut_13_1 (
    .O(x13_y1),
    .I0(x11_y5),
    .I1(x10_y3),
    .I2(1'b0),
    .I3(x10_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110110100110)
) lut_14_1 (
    .O(x14_y1),
    .I0(x11_y5),
    .I1(x12_y4),
    .I2(x12_y0),
    .I3(x12_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110010000110)
) lut_15_1 (
    .O(x15_y1),
    .I0(1'b0),
    .I1(x12_y2),
    .I2(x12_y2),
    .I3(x13_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011110001000)
) lut_16_1 (
    .O(x16_y1),
    .I0(x13_y0),
    .I1(x14_y5),
    .I2(x14_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010100100101)
) lut_17_1 (
    .O(x17_y1),
    .I0(x15_y6),
    .I1(x14_y6),
    .I2(x14_y2),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100101110101)
) lut_18_1 (
    .O(x18_y1),
    .I0(x15_y4),
    .I1(x16_y0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100011111010)
) lut_19_1 (
    .O(x19_y1),
    .I0(x16_y1),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x16_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001010100011)
) lut_20_1 (
    .O(x20_y1),
    .I0(x18_y6),
    .I1(x17_y1),
    .I2(x18_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110010000011)
) lut_21_1 (
    .O(x21_y1),
    .I0(x19_y5),
    .I1(x19_y0),
    .I2(x19_y0),
    .I3(x18_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110111110010)
) lut_22_1 (
    .O(x22_y1),
    .I0(x20_y3),
    .I1(1'b0),
    .I2(x20_y0),
    .I3(x19_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001001111010)
) lut_23_1 (
    .O(x23_y1),
    .I0(1'b0),
    .I1(x21_y4),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110001011101)
) lut_24_1 (
    .O(x24_y1),
    .I0(x22_y2),
    .I1(x22_y6),
    .I2(x22_y2),
    .I3(x22_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101000001111)
) lut_25_1 (
    .O(x25_y1),
    .I0(x23_y0),
    .I1(x22_y2),
    .I2(x23_y1),
    .I3(x23_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101111101100)
) lut_26_1 (
    .O(x26_y1),
    .I0(x24_y5),
    .I1(x24_y1),
    .I2(x24_y2),
    .I3(x23_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110000000010)
) lut_27_1 (
    .O(x27_y1),
    .I0(x24_y3),
    .I1(1'b0),
    .I2(x24_y5),
    .I3(x24_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011011000111)
) lut_28_1 (
    .O(x28_y1),
    .I0(x26_y0),
    .I1(x25_y3),
    .I2(x26_y6),
    .I3(x26_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010000000000)
) lut_29_1 (
    .O(x29_y1),
    .I0(x27_y2),
    .I1(x27_y2),
    .I2(x27_y3),
    .I3(x27_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110100001000)
) lut_30_1 (
    .O(x30_y1),
    .I0(x28_y4),
    .I1(1'b0),
    .I2(x27_y6),
    .I3(x27_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001010110010)
) lut_31_1 (
    .O(x31_y1),
    .I0(x28_y4),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111111000011)
) lut_32_1 (
    .O(x32_y1),
    .I0(x29_y3),
    .I1(1'b0),
    .I2(x30_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001011101000)
) lut_33_1 (
    .O(x33_y1),
    .I0(x30_y0),
    .I1(x30_y0),
    .I2(x30_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110011100011)
) lut_34_1 (
    .O(x34_y1),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x32_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111111010011)
) lut_35_1 (
    .O(x35_y1),
    .I0(x32_y0),
    .I1(x32_y1),
    .I2(1'b0),
    .I3(x32_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100101111011)
) lut_36_1 (
    .O(x36_y1),
    .I0(x34_y0),
    .I1(x34_y5),
    .I2(x34_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000101001110)
) lut_37_1 (
    .O(x37_y1),
    .I0(1'b0),
    .I1(x34_y1),
    .I2(x34_y5),
    .I3(x35_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010111111110)
) lut_38_1 (
    .O(x38_y1),
    .I0(x35_y6),
    .I1(1'b0),
    .I2(x35_y6),
    .I3(x35_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011101011110)
) lut_39_1 (
    .O(x39_y1),
    .I0(x36_y0),
    .I1(x37_y5),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000101000101)
) lut_40_1 (
    .O(x40_y1),
    .I0(x38_y0),
    .I1(x37_y4),
    .I2(x38_y6),
    .I3(x37_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100100110110)
) lut_41_1 (
    .O(x41_y1),
    .I0(x38_y2),
    .I1(x39_y0),
    .I2(1'b0),
    .I3(x39_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010000110110)
) lut_42_1 (
    .O(x42_y1),
    .I0(x39_y0),
    .I1(x39_y0),
    .I2(1'b0),
    .I3(x40_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011000111000)
) lut_43_1 (
    .O(x43_y1),
    .I0(x41_y0),
    .I1(x40_y0),
    .I2(1'b0),
    .I3(x41_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001101111111)
) lut_44_1 (
    .O(x44_y1),
    .I0(x41_y0),
    .I1(x42_y0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100110111001)
) lut_45_1 (
    .O(x45_y1),
    .I0(1'b0),
    .I1(x42_y1),
    .I2(x42_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001110111011)
) lut_46_1 (
    .O(x46_y1),
    .I0(x44_y3),
    .I1(x43_y2),
    .I2(x44_y1),
    .I3(x44_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000101111100)
) lut_47_1 (
    .O(x47_y1),
    .I0(x45_y5),
    .I1(x45_y2),
    .I2(x45_y2),
    .I3(x44_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101001100110)
) lut_48_1 (
    .O(x48_y1),
    .I0(x45_y0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x45_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010100001000)
) lut_49_1 (
    .O(x49_y1),
    .I0(1'b0),
    .I1(x47_y6),
    .I2(1'b0),
    .I3(x46_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000110100100)
) lut_50_1 (
    .O(x50_y1),
    .I0(1'b0),
    .I1(x47_y4),
    .I2(x47_y0),
    .I3(x48_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100101001111)
) lut_51_1 (
    .O(x51_y1),
    .I0(x49_y4),
    .I1(x49_y5),
    .I2(x49_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101101101001)
) lut_52_1 (
    .O(x52_y1),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100110110000)
) lut_53_1 (
    .O(x53_y1),
    .I0(x51_y5),
    .I1(1'b0),
    .I2(x50_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100111100011)
) lut_54_1 (
    .O(x54_y1),
    .I0(x52_y2),
    .I1(x52_y0),
    .I2(x52_y6),
    .I3(x52_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001110110111)
) lut_55_1 (
    .O(x55_y1),
    .I0(x52_y4),
    .I1(x53_y6),
    .I2(x52_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001000000111)
) lut_56_1 (
    .O(x56_y1),
    .I0(x53_y2),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x54_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010111010111)
) lut_57_1 (
    .O(x57_y1),
    .I0(1'b0),
    .I1(x55_y0),
    .I2(x55_y1),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000101001110)
) lut_58_1 (
    .O(x58_y1),
    .I0(x55_y3),
    .I1(x56_y5),
    .I2(x55_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100011010001)
) lut_59_1 (
    .O(x59_y1),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x56_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011110101010)
) lut_60_1 (
    .O(x60_y1),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x58_y0),
    .I3(x57_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100111101010)
) lut_61_1 (
    .O(x61_y1),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x58_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110001110011)
) lut_62_1 (
    .O(x62_y1),
    .I0(x60_y0),
    .I1(x59_y5),
    .I2(1'b0),
    .I3(x60_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010100011001)
) lut_0_2 (
    .O(x0_y2),
    .I0(in2),
    .I1(in6),
    .I2(in7),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010110011111)
) lut_1_2 (
    .O(x1_y2),
    .I0(in6),
    .I1(in7),
    .I2(1'b0),
    .I3(in5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000110110110)
) lut_2_2 (
    .O(x2_y2),
    .I0(1'b0),
    .I1(in7),
    .I2(1'b0),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111000100101)
) lut_3_2 (
    .O(x3_y2),
    .I0(in0),
    .I1(x1_y6),
    .I2(in4),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100111100010)
) lut_4_2 (
    .O(x4_y2),
    .I0(x2_y5),
    .I1(x2_y0),
    .I2(x2_y0),
    .I3(x1_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100101100011)
) lut_5_2 (
    .O(x5_y2),
    .I0(x3_y0),
    .I1(1'b0),
    .I2(x3_y2),
    .I3(x2_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111000001001)
) lut_6_2 (
    .O(x6_y2),
    .I0(x4_y0),
    .I1(x3_y3),
    .I2(x4_y6),
    .I3(x3_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000100100010)
) lut_7_2 (
    .O(x7_y2),
    .I0(x4_y3),
    .I1(x5_y4),
    .I2(x4_y7),
    .I3(x5_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110011100110)
) lut_8_2 (
    .O(x8_y2),
    .I0(x6_y4),
    .I1(x6_y7),
    .I2(x5_y0),
    .I3(x6_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101000101101)
) lut_9_2 (
    .O(x9_y2),
    .I0(x6_y3),
    .I1(x7_y0),
    .I2(x5_y0),
    .I3(x6_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110001111110)
) lut_10_2 (
    .O(x10_y2),
    .I0(x8_y1),
    .I1(x8_y0),
    .I2(1'b0),
    .I3(x8_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010111101011)
) lut_11_2 (
    .O(x11_y2),
    .I0(1'b0),
    .I1(x9_y0),
    .I2(x8_y7),
    .I3(x8_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010111000010)
) lut_12_2 (
    .O(x12_y2),
    .I0(1'b0),
    .I1(x10_y4),
    .I2(x9_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110100100110)
) lut_13_2 (
    .O(x13_y2),
    .I0(1'b0),
    .I1(x11_y0),
    .I2(x11_y0),
    .I3(x11_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011111010011)
) lut_14_2 (
    .O(x14_y2),
    .I0(1'b0),
    .I1(x11_y4),
    .I2(x11_y4),
    .I3(x12_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100101101001)
) lut_15_2 (
    .O(x15_y2),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x12_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011010000101)
) lut_16_2 (
    .O(x16_y2),
    .I0(x13_y3),
    .I1(x14_y0),
    .I2(x14_y5),
    .I3(x13_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110100110001)
) lut_17_2 (
    .O(x17_y2),
    .I0(x14_y0),
    .I1(1'b0),
    .I2(x14_y0),
    .I3(x15_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110101000010)
) lut_18_2 (
    .O(x18_y2),
    .I0(1'b0),
    .I1(x15_y7),
    .I2(x15_y0),
    .I3(x15_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101100100010)
) lut_19_2 (
    .O(x19_y2),
    .I0(x16_y1),
    .I1(1'b0),
    .I2(x16_y4),
    .I3(x16_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011000001011)
) lut_20_2 (
    .O(x20_y2),
    .I0(x18_y5),
    .I1(x18_y0),
    .I2(x17_y0),
    .I3(x17_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000111111111)
) lut_21_2 (
    .O(x21_y2),
    .I0(x19_y5),
    .I1(1'b0),
    .I2(x19_y1),
    .I3(x18_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100110010100)
) lut_22_2 (
    .O(x22_y2),
    .I0(x20_y0),
    .I1(x20_y0),
    .I2(1'b0),
    .I3(x19_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000010010110)
) lut_23_2 (
    .O(x23_y2),
    .I0(x20_y0),
    .I1(x20_y4),
    .I2(x20_y5),
    .I3(x21_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001011000011)
) lut_24_2 (
    .O(x24_y2),
    .I0(x22_y0),
    .I1(x22_y7),
    .I2(x21_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100010001000)
) lut_25_2 (
    .O(x25_y2),
    .I0(x23_y6),
    .I1(1'b0),
    .I2(x22_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011001111110)
) lut_26_2 (
    .O(x26_y2),
    .I0(x23_y0),
    .I1(x23_y6),
    .I2(x24_y6),
    .I3(x24_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111100001011)
) lut_27_2 (
    .O(x27_y2),
    .I0(x24_y0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111101111110)
) lut_28_2 (
    .O(x28_y2),
    .I0(x26_y0),
    .I1(x25_y0),
    .I2(x25_y0),
    .I3(x25_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000011101011)
) lut_29_2 (
    .O(x29_y2),
    .I0(x27_y6),
    .I1(x26_y5),
    .I2(x27_y1),
    .I3(x26_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100111110001)
) lut_30_2 (
    .O(x30_y2),
    .I0(x27_y7),
    .I1(x27_y4),
    .I2(x27_y5),
    .I3(x28_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111100001010)
) lut_31_2 (
    .O(x31_y2),
    .I0(x29_y0),
    .I1(1'b0),
    .I2(x28_y0),
    .I3(x29_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001100111110)
) lut_32_2 (
    .O(x32_y2),
    .I0(x29_y4),
    .I1(x29_y1),
    .I2(1'b0),
    .I3(x29_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000101110110)
) lut_33_2 (
    .O(x33_y2),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x31_y2),
    .I3(x30_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111011001110)
) lut_34_2 (
    .O(x34_y2),
    .I0(x32_y2),
    .I1(x32_y2),
    .I2(1'b0),
    .I3(x32_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110101111001)
) lut_35_2 (
    .O(x35_y2),
    .I0(x32_y2),
    .I1(x33_y1),
    .I2(x33_y2),
    .I3(x32_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011011011011)
) lut_36_2 (
    .O(x36_y2),
    .I0(x34_y5),
    .I1(x34_y4),
    .I2(1'b0),
    .I3(x34_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010100001111)
) lut_37_2 (
    .O(x37_y2),
    .I0(1'b0),
    .I1(x34_y2),
    .I2(1'b0),
    .I3(x34_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111000110010)
) lut_38_2 (
    .O(x38_y2),
    .I0(x36_y1),
    .I1(x36_y1),
    .I2(1'b0),
    .I3(x36_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001101110101)
) lut_39_2 (
    .O(x39_y2),
    .I0(x37_y0),
    .I1(x36_y0),
    .I2(1'b0),
    .I3(x36_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111100100110)
) lut_40_2 (
    .O(x40_y2),
    .I0(x37_y5),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x37_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001000111111)
) lut_41_2 (
    .O(x41_y2),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x39_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110100100011)
) lut_42_2 (
    .O(x42_y2),
    .I0(x39_y0),
    .I1(x40_y0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100011011001)
) lut_43_2 (
    .O(x43_y2),
    .I0(1'b0),
    .I1(x40_y0),
    .I2(x40_y0),
    .I3(x40_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010001100101)
) lut_44_2 (
    .O(x44_y2),
    .I0(x42_y2),
    .I1(x41_y7),
    .I2(1'b0),
    .I3(x41_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100011100010)
) lut_45_2 (
    .O(x45_y2),
    .I0(1'b0),
    .I1(x43_y0),
    .I2(x43_y2),
    .I3(x42_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001101010001)
) lut_46_2 (
    .O(x46_y2),
    .I0(x43_y0),
    .I1(x44_y2),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001100100111)
) lut_47_2 (
    .O(x47_y2),
    .I0(x44_y0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x45_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000110101100)
) lut_48_2 (
    .O(x48_y2),
    .I0(x45_y3),
    .I1(x45_y0),
    .I2(x45_y6),
    .I3(x46_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001110100111)
) lut_49_2 (
    .O(x49_y2),
    .I0(x47_y6),
    .I1(x47_y2),
    .I2(x46_y4),
    .I3(x46_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111101010001)
) lut_50_2 (
    .O(x50_y2),
    .I0(1'b0),
    .I1(x48_y3),
    .I2(x48_y0),
    .I3(x47_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010110110001)
) lut_51_2 (
    .O(x51_y2),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x49_y0),
    .I3(x49_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001100110101)
) lut_52_2 (
    .O(x52_y2),
    .I0(x49_y0),
    .I1(x49_y4),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001011101011)
) lut_53_2 (
    .O(x53_y2),
    .I0(x50_y1),
    .I1(x51_y5),
    .I2(x50_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111010110101)
) lut_54_2 (
    .O(x54_y2),
    .I0(x51_y6),
    .I1(x51_y1),
    .I2(x51_y0),
    .I3(x52_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011110110001)
) lut_55_2 (
    .O(x55_y2),
    .I0(x53_y7),
    .I1(x52_y0),
    .I2(x52_y1),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011010100110)
) lut_56_2 (
    .O(x56_y2),
    .I0(x54_y4),
    .I1(1'b0),
    .I2(x54_y7),
    .I3(x54_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000010111001)
) lut_57_2 (
    .O(x57_y2),
    .I0(1'b0),
    .I1(x55_y7),
    .I2(x55_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111001001100)
) lut_58_2 (
    .O(x58_y2),
    .I0(x56_y1),
    .I1(x55_y6),
    .I2(x55_y3),
    .I3(x56_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011111111100)
) lut_59_2 (
    .O(x59_y2),
    .I0(x57_y3),
    .I1(x56_y0),
    .I2(x56_y0),
    .I3(x56_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000001111111)
) lut_60_2 (
    .O(x60_y2),
    .I0(x57_y0),
    .I1(x58_y6),
    .I2(1'b0),
    .I3(x57_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000001000010)
) lut_61_2 (
    .O(x61_y2),
    .I0(x58_y1),
    .I1(x59_y0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100110010001)
) lut_62_2 (
    .O(x62_y2),
    .I0(x60_y0),
    .I1(x60_y0),
    .I2(1'b0),
    .I3(x59_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100000000000)
) lut_0_3 (
    .O(x0_y3),
    .I0(in6),
    .I1(1'b0),
    .I2(in1),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111010010100)
) lut_1_3 (
    .O(x1_y3),
    .I0(1'b0),
    .I1(in7),
    .I2(in3),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100101010101)
) lut_2_3 (
    .O(x2_y3),
    .I0(1'b0),
    .I1(in6),
    .I2(1'b0),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010000101110)
) lut_3_3 (
    .O(x3_y3),
    .I0(1'b0),
    .I1(in6),
    .I2(in0),
    .I3(x1_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111101101100)
) lut_4_3 (
    .O(x4_y3),
    .I0(x2_y4),
    .I1(x1_y6),
    .I2(x1_y7),
    .I3(x1_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011110010011)
) lut_5_3 (
    .O(x5_y3),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x3_y8),
    .I3(x2_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001100001010)
) lut_6_3 (
    .O(x6_y3),
    .I0(x4_y0),
    .I1(x3_y0),
    .I2(x3_y1),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110010101101)
) lut_7_3 (
    .O(x7_y3),
    .I0(x4_y3),
    .I1(x5_y8),
    .I2(x5_y4),
    .I3(x5_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000100110111)
) lut_8_3 (
    .O(x8_y3),
    .I0(x5_y2),
    .I1(x5_y0),
    .I2(x6_y3),
    .I3(x6_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010111110010)
) lut_9_3 (
    .O(x9_y3),
    .I0(x7_y4),
    .I1(1'b0),
    .I2(x6_y3),
    .I3(x6_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000110101010)
) lut_10_3 (
    .O(x10_y3),
    .I0(x8_y0),
    .I1(x8_y4),
    .I2(x8_y0),
    .I3(x7_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101100011110)
) lut_11_3 (
    .O(x11_y3),
    .I0(x9_y5),
    .I1(x9_y6),
    .I2(x9_y0),
    .I3(x9_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001001010001)
) lut_12_3 (
    .O(x12_y3),
    .I0(x10_y1),
    .I1(x9_y1),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110100000101)
) lut_13_3 (
    .O(x13_y3),
    .I0(x10_y0),
    .I1(x11_y3),
    .I2(x10_y3),
    .I3(x11_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111111110001)
) lut_14_3 (
    .O(x14_y3),
    .I0(x12_y0),
    .I1(x11_y4),
    .I2(1'b0),
    .I3(x11_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000001111100)
) lut_15_3 (
    .O(x15_y3),
    .I0(1'b0),
    .I1(x13_y4),
    .I2(x12_y7),
    .I3(x13_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101001001010)
) lut_16_3 (
    .O(x16_y3),
    .I0(1'b0),
    .I1(x14_y2),
    .I2(x14_y2),
    .I3(x14_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000001000011)
) lut_17_3 (
    .O(x17_y3),
    .I0(x15_y1),
    .I1(1'b0),
    .I2(x15_y1),
    .I3(x15_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010000010100)
) lut_18_3 (
    .O(x18_y3),
    .I0(x15_y0),
    .I1(x16_y2),
    .I2(x15_y2),
    .I3(x16_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000001001010)
) lut_19_3 (
    .O(x19_y3),
    .I0(1'b0),
    .I1(x17_y2),
    .I2(1'b0),
    .I3(x17_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100000001011)
) lut_20_3 (
    .O(x20_y3),
    .I0(x18_y6),
    .I1(x18_y6),
    .I2(x18_y2),
    .I3(x17_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111110010111)
) lut_21_3 (
    .O(x21_y3),
    .I0(x18_y5),
    .I1(x18_y8),
    .I2(x18_y4),
    .I3(x19_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110100100110)
) lut_22_3 (
    .O(x22_y3),
    .I0(x19_y8),
    .I1(x19_y0),
    .I2(1'b0),
    .I3(x20_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011001101100)
) lut_23_3 (
    .O(x23_y3),
    .I0(1'b0),
    .I1(x21_y3),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100001001011)
) lut_24_3 (
    .O(x24_y3),
    .I0(x21_y0),
    .I1(x22_y1),
    .I2(x21_y4),
    .I3(x22_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101110011110)
) lut_25_3 (
    .O(x25_y3),
    .I0(x22_y6),
    .I1(x23_y2),
    .I2(x22_y0),
    .I3(x22_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101110110110)
) lut_26_3 (
    .O(x26_y3),
    .I0(x24_y0),
    .I1(x23_y1),
    .I2(x23_y0),
    .I3(x24_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101000011101)
) lut_27_3 (
    .O(x27_y3),
    .I0(1'b0),
    .I1(x24_y0),
    .I2(x24_y1),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110111011110)
) lut_28_3 (
    .O(x28_y3),
    .I0(1'b0),
    .I1(x26_y8),
    .I2(x26_y6),
    .I3(x25_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000111011000)
) lut_29_3 (
    .O(x29_y3),
    .I0(x27_y8),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x27_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111101010110)
) lut_30_3 (
    .O(x30_y3),
    .I0(x28_y0),
    .I1(x28_y1),
    .I2(x27_y1),
    .I3(x28_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010101010100)
) lut_31_3 (
    .O(x31_y3),
    .I0(x29_y2),
    .I1(x29_y7),
    .I2(x29_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010100100101)
) lut_32_3 (
    .O(x32_y3),
    .I0(x30_y0),
    .I1(x29_y7),
    .I2(x30_y1),
    .I3(x30_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110011100000)
) lut_33_3 (
    .O(x33_y3),
    .I0(x31_y6),
    .I1(x31_y8),
    .I2(x30_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010101001000)
) lut_34_3 (
    .O(x34_y3),
    .I0(x32_y7),
    .I1(x32_y0),
    .I2(x32_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110100111011)
) lut_35_3 (
    .O(x35_y3),
    .I0(x33_y8),
    .I1(x32_y0),
    .I2(1'b0),
    .I3(x33_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110101111010)
) lut_36_3 (
    .O(x36_y3),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x33_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111000100101)
) lut_37_3 (
    .O(x37_y3),
    .I0(x35_y8),
    .I1(x34_y0),
    .I2(x35_y0),
    .I3(x34_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111110110011)
) lut_38_3 (
    .O(x38_y3),
    .I0(1'b0),
    .I1(x36_y0),
    .I2(x36_y4),
    .I3(x35_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111100110110)
) lut_39_3 (
    .O(x39_y3),
    .I0(x37_y6),
    .I1(1'b0),
    .I2(x37_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010000010011)
) lut_40_3 (
    .O(x40_y3),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x37_y6),
    .I3(x38_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100001000011)
) lut_41_3 (
    .O(x41_y3),
    .I0(x39_y8),
    .I1(x38_y5),
    .I2(x38_y3),
    .I3(x38_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010100101000)
) lut_42_3 (
    .O(x42_y3),
    .I0(x40_y1),
    .I1(x39_y2),
    .I2(x39_y4),
    .I3(x39_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101101111011)
) lut_43_3 (
    .O(x43_y3),
    .I0(x41_y6),
    .I1(x41_y0),
    .I2(x41_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100000100111)
) lut_44_3 (
    .O(x44_y3),
    .I0(x42_y2),
    .I1(x42_y6),
    .I2(1'b0),
    .I3(x42_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111001011100)
) lut_45_3 (
    .O(x45_y3),
    .I0(x43_y8),
    .I1(x42_y6),
    .I2(1'b0),
    .I3(x42_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001010111001)
) lut_46_3 (
    .O(x46_y3),
    .I0(x43_y5),
    .I1(x43_y0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010001001110)
) lut_47_3 (
    .O(x47_y3),
    .I0(x45_y8),
    .I1(1'b0),
    .I2(x44_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111010000001)
) lut_48_3 (
    .O(x48_y3),
    .I0(x45_y0),
    .I1(1'b0),
    .I2(x46_y0),
    .I3(x46_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111101011100)
) lut_49_3 (
    .O(x49_y3),
    .I0(x47_y3),
    .I1(x46_y5),
    .I2(x47_y0),
    .I3(x46_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111111001111)
) lut_50_3 (
    .O(x50_y3),
    .I0(x47_y1),
    .I1(x48_y6),
    .I2(x48_y0),
    .I3(x47_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101001000100)
) lut_51_3 (
    .O(x51_y3),
    .I0(x48_y3),
    .I1(x49_y1),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001011111000)
) lut_52_3 (
    .O(x52_y3),
    .I0(x49_y7),
    .I1(x49_y6),
    .I2(x49_y7),
    .I3(x49_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000111011001)
) lut_53_3 (
    .O(x53_y3),
    .I0(x50_y8),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010000100101)
) lut_54_3 (
    .O(x54_y3),
    .I0(x52_y7),
    .I1(1'b0),
    .I2(x52_y0),
    .I3(x51_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110011111000)
) lut_55_3 (
    .O(x55_y3),
    .I0(x53_y8),
    .I1(1'b0),
    .I2(x53_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110000001000)
) lut_56_3 (
    .O(x56_y3),
    .I0(1'b0),
    .I1(x54_y5),
    .I2(x54_y0),
    .I3(x53_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011110000001)
) lut_57_3 (
    .O(x57_y3),
    .I0(x55_y7),
    .I1(x55_y0),
    .I2(1'b0),
    .I3(x55_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110010011001)
) lut_58_3 (
    .O(x58_y3),
    .I0(x55_y0),
    .I1(x56_y0),
    .I2(x56_y8),
    .I3(x56_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101110001010)
) lut_59_3 (
    .O(x59_y3),
    .I0(x57_y1),
    .I1(x57_y0),
    .I2(x57_y7),
    .I3(x57_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110110010011)
) lut_60_3 (
    .O(x60_y3),
    .I0(x58_y6),
    .I1(x57_y1),
    .I2(x58_y0),
    .I3(x57_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010101010000)
) lut_61_3 (
    .O(x61_y3),
    .I0(x58_y1),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x59_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011110101010)
) lut_62_3 (
    .O(x62_y3),
    .I0(x59_y7),
    .I1(x60_y0),
    .I2(x60_y1),
    .I3(x60_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100000000011)
) lut_0_4 (
    .O(x0_y4),
    .I0(in3),
    .I1(1'b0),
    .I2(in0),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010010110001)
) lut_1_4 (
    .O(x1_y4),
    .I0(in9),
    .I1(in8),
    .I2(in7),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100111011000)
) lut_2_4 (
    .O(x2_y4),
    .I0(1'b0),
    .I1(1'b0),
    .I2(in3),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111101100111)
) lut_3_4 (
    .O(x3_y4),
    .I0(x1_y4),
    .I1(1'b0),
    .I2(in1),
    .I3(x1_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111000101100)
) lut_4_4 (
    .O(x4_y4),
    .I0(x1_y9),
    .I1(x2_y4),
    .I2(x2_y1),
    .I3(x2_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101000001110)
) lut_5_4 (
    .O(x5_y4),
    .I0(1'b0),
    .I1(x2_y8),
    .I2(x3_y6),
    .I3(x3_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001101101000)
) lut_6_4 (
    .O(x6_y4),
    .I0(x4_y0),
    .I1(x3_y3),
    .I2(x4_y3),
    .I3(x3_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011000101110)
) lut_7_4 (
    .O(x7_y4),
    .I0(x4_y3),
    .I1(x5_y5),
    .I2(x5_y5),
    .I3(x4_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100000001110)
) lut_8_4 (
    .O(x8_y4),
    .I0(x6_y5),
    .I1(x6_y1),
    .I2(x5_y5),
    .I3(x6_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010101011110)
) lut_9_4 (
    .O(x9_y4),
    .I0(1'b0),
    .I1(x7_y2),
    .I2(x5_y5),
    .I3(x6_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000010110111)
) lut_10_4 (
    .O(x10_y4),
    .I0(x7_y0),
    .I1(x7_y7),
    .I2(x8_y2),
    .I3(x7_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110010111100)
) lut_11_4 (
    .O(x11_y4),
    .I0(1'b0),
    .I1(x8_y2),
    .I2(1'b0),
    .I3(x9_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101000000000)
) lut_12_4 (
    .O(x12_y4),
    .I0(x10_y4),
    .I1(1'b0),
    .I2(x10_y0),
    .I3(x9_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110100010000)
) lut_13_4 (
    .O(x13_y4),
    .I0(x10_y7),
    .I1(x11_y9),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010100100100)
) lut_14_4 (
    .O(x14_y4),
    .I0(x11_y2),
    .I1(1'b0),
    .I2(x11_y1),
    .I3(x12_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010111110011)
) lut_15_4 (
    .O(x15_y4),
    .I0(x12_y1),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001010001100)
) lut_16_4 (
    .O(x16_y4),
    .I0(1'b0),
    .I1(x14_y0),
    .I2(x14_y2),
    .I3(x14_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010001010101)
) lut_17_4 (
    .O(x17_y4),
    .I0(x15_y2),
    .I1(x14_y0),
    .I2(x15_y6),
    .I3(x15_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011010101001)
) lut_18_4 (
    .O(x18_y4),
    .I0(1'b0),
    .I1(x16_y3),
    .I2(1'b0),
    .I3(x15_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111100001000)
) lut_19_4 (
    .O(x19_y4),
    .I0(x16_y2),
    .I1(x16_y6),
    .I2(x16_y7),
    .I3(x16_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010111100011)
) lut_20_4 (
    .O(x20_y4),
    .I0(x18_y4),
    .I1(1'b0),
    .I2(x17_y2),
    .I3(x18_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010100110111)
) lut_21_4 (
    .O(x21_y4),
    .I0(x19_y7),
    .I1(x18_y2),
    .I2(1'b0),
    .I3(x18_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110000111010)
) lut_22_4 (
    .O(x22_y4),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100110011111)
) lut_23_4 (
    .O(x23_y4),
    .I0(x21_y8),
    .I1(1'b0),
    .I2(x20_y3),
    .I3(x20_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111110101100)
) lut_24_4 (
    .O(x24_y4),
    .I0(1'b0),
    .I1(x21_y4),
    .I2(1'b0),
    .I3(x22_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100001000101)
) lut_25_4 (
    .O(x25_y4),
    .I0(x23_y1),
    .I1(x22_y2),
    .I2(x22_y7),
    .I3(x22_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010000011001)
) lut_26_4 (
    .O(x26_y4),
    .I0(1'b0),
    .I1(x23_y5),
    .I2(x23_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101111110111)
) lut_27_4 (
    .O(x27_y4),
    .I0(x25_y8),
    .I1(x24_y7),
    .I2(x24_y7),
    .I3(x25_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000001010100)
) lut_28_4 (
    .O(x28_y4),
    .I0(1'b0),
    .I1(x26_y5),
    .I2(x25_y4),
    .I3(x26_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100100011110)
) lut_29_4 (
    .O(x29_y4),
    .I0(1'b0),
    .I1(x26_y7),
    .I2(x26_y0),
    .I3(x26_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001010010010)
) lut_30_4 (
    .O(x30_y4),
    .I0(x27_y7),
    .I1(x28_y7),
    .I2(x28_y8),
    .I3(x27_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011010010110)
) lut_31_4 (
    .O(x31_y4),
    .I0(x29_y0),
    .I1(x29_y4),
    .I2(x28_y9),
    .I3(x29_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010101100100)
) lut_32_4 (
    .O(x32_y4),
    .I0(1'b0),
    .I1(x29_y5),
    .I2(x30_y7),
    .I3(x29_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001110010101)
) lut_33_4 (
    .O(x33_y4),
    .I0(x31_y0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x31_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101100010111)
) lut_34_4 (
    .O(x34_y4),
    .I0(x31_y1),
    .I1(x32_y8),
    .I2(x31_y9),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001010001110)
) lut_35_4 (
    .O(x35_y4),
    .I0(x32_y0),
    .I1(x32_y0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100011001001)
) lut_36_4 (
    .O(x36_y4),
    .I0(x34_y3),
    .I1(1'b0),
    .I2(x34_y7),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110000110000)
) lut_37_4 (
    .O(x37_y4),
    .I0(x35_y2),
    .I1(x35_y5),
    .I2(x34_y1),
    .I3(x35_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001000001010)
) lut_38_4 (
    .O(x38_y4),
    .I0(x36_y3),
    .I1(x35_y4),
    .I2(x36_y6),
    .I3(x35_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011000010100)
) lut_39_4 (
    .O(x39_y4),
    .I0(x37_y7),
    .I1(x36_y3),
    .I2(x37_y0),
    .I3(x37_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000110010110)
) lut_40_4 (
    .O(x40_y4),
    .I0(x38_y0),
    .I1(x38_y0),
    .I2(x37_y8),
    .I3(x37_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110111100111)
) lut_41_4 (
    .O(x41_y4),
    .I0(x39_y3),
    .I1(x39_y2),
    .I2(x38_y1),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011010010110)
) lut_42_4 (
    .O(x42_y4),
    .I0(x39_y7),
    .I1(x40_y5),
    .I2(x40_y4),
    .I3(x40_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001100101010)
) lut_43_4 (
    .O(x43_y4),
    .I0(x41_y0),
    .I1(x40_y0),
    .I2(1'b0),
    .I3(x40_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100101001110)
) lut_44_4 (
    .O(x44_y4),
    .I0(x41_y8),
    .I1(x42_y6),
    .I2(x42_y7),
    .I3(x41_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011111000001)
) lut_45_4 (
    .O(x45_y4),
    .I0(x42_y0),
    .I1(1'b0),
    .I2(x42_y8),
    .I3(x42_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001101110110)
) lut_46_4 (
    .O(x46_y4),
    .I0(1'b0),
    .I1(x44_y4),
    .I2(1'b0),
    .I3(x44_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010010111110)
) lut_47_4 (
    .O(x47_y4),
    .I0(x44_y8),
    .I1(x44_y2),
    .I2(x44_y5),
    .I3(x44_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001101011100)
) lut_48_4 (
    .O(x48_y4),
    .I0(x45_y0),
    .I1(x45_y5),
    .I2(1'b0),
    .I3(x46_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100101110111)
) lut_49_4 (
    .O(x49_y4),
    .I0(x47_y1),
    .I1(x46_y8),
    .I2(x46_y7),
    .I3(x46_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110110001001)
) lut_50_4 (
    .O(x50_y4),
    .I0(x48_y6),
    .I1(1'b0),
    .I2(x47_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011001011001)
) lut_51_4 (
    .O(x51_y4),
    .I0(x49_y4),
    .I1(x48_y0),
    .I2(x48_y9),
    .I3(x48_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110000001011)
) lut_52_4 (
    .O(x52_y4),
    .I0(x49_y2),
    .I1(x49_y2),
    .I2(x50_y2),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111000001000)
) lut_53_4 (
    .O(x53_y4),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x51_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110111000100)
) lut_54_4 (
    .O(x54_y4),
    .I0(x51_y6),
    .I1(1'b0),
    .I2(x52_y8),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101101101010)
) lut_55_4 (
    .O(x55_y4),
    .I0(x53_y7),
    .I1(1'b0),
    .I2(x53_y7),
    .I3(x53_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011011001000)
) lut_56_4 (
    .O(x56_y4),
    .I0(x54_y2),
    .I1(1'b0),
    .I2(x54_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111110000111)
) lut_57_4 (
    .O(x57_y4),
    .I0(x54_y0),
    .I1(x55_y7),
    .I2(1'b0),
    .I3(x55_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000100111010)
) lut_58_4 (
    .O(x58_y4),
    .I0(x56_y5),
    .I1(1'b0),
    .I2(x56_y0),
    .I3(x55_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111110110101)
) lut_59_4 (
    .O(x59_y4),
    .I0(x57_y2),
    .I1(x56_y0),
    .I2(1'b0),
    .I3(x56_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011001110010)
) lut_60_4 (
    .O(x60_y4),
    .I0(x58_y6),
    .I1(x57_y7),
    .I2(x57_y9),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001010110000)
) lut_61_4 (
    .O(x61_y4),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x58_y0),
    .I3(x58_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111110000100)
) lut_62_4 (
    .O(x62_y4),
    .I0(1'b0),
    .I1(x60_y1),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101001001011)
) lut_0_5 (
    .O(x0_y5),
    .I0(in8),
    .I1(in4),
    .I2(in4),
    .I3(in7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100110001001)
) lut_1_5 (
    .O(x1_y5),
    .I0(in1),
    .I1(in3),
    .I2(in4),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100101100100)
) lut_2_5 (
    .O(x2_y5),
    .I0(in7),
    .I1(1'b0),
    .I2(in0),
    .I3(in9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000110110010)
) lut_3_5 (
    .O(x3_y5),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x1_y9),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011101110101)
) lut_4_5 (
    .O(x4_y5),
    .I0(x2_y0),
    .I1(x1_y10),
    .I2(x1_y9),
    .I3(x1_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101101001001)
) lut_5_5 (
    .O(x5_y5),
    .I0(x2_y3),
    .I1(x3_y9),
    .I2(x2_y3),
    .I3(x3_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011000001011)
) lut_6_5 (
    .O(x6_y5),
    .I0(x3_y6),
    .I1(x4_y10),
    .I2(1'b0),
    .I3(x4_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100111010110)
) lut_7_5 (
    .O(x7_y5),
    .I0(1'b0),
    .I1(x4_y9),
    .I2(x5_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100011101111)
) lut_8_5 (
    .O(x8_y5),
    .I0(x5_y5),
    .I1(x6_y9),
    .I2(1'b0),
    .I3(x5_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000101101001)
) lut_9_5 (
    .O(x9_y5),
    .I0(x6_y0),
    .I1(x6_y4),
    .I2(1'b0),
    .I3(x5_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000001000100)
) lut_10_5 (
    .O(x10_y5),
    .I0(1'b0),
    .I1(x7_y0),
    .I2(x7_y4),
    .I3(x7_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000110010001)
) lut_11_5 (
    .O(x11_y5),
    .I0(x9_y6),
    .I1(x8_y5),
    .I2(x8_y7),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101010110101)
) lut_12_5 (
    .O(x12_y5),
    .I0(x9_y4),
    .I1(x10_y10),
    .I2(x10_y10),
    .I3(x10_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101010111000)
) lut_13_5 (
    .O(x13_y5),
    .I0(1'b0),
    .I1(x10_y7),
    .I2(1'b0),
    .I3(x10_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010100000110)
) lut_14_5 (
    .O(x14_y5),
    .I0(x12_y7),
    .I1(x12_y10),
    .I2(x12_y2),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101000010011)
) lut_15_5 (
    .O(x15_y5),
    .I0(x12_y3),
    .I1(x12_y3),
    .I2(x12_y1),
    .I3(x13_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111110010111)
) lut_16_5 (
    .O(x16_y5),
    .I0(x13_y1),
    .I1(x14_y9),
    .I2(x13_y0),
    .I3(x14_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001110111100)
) lut_17_5 (
    .O(x17_y5),
    .I0(1'b0),
    .I1(x14_y0),
    .I2(x14_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100111100011)
) lut_18_5 (
    .O(x18_y5),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x15_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110111100001)
) lut_19_5 (
    .O(x19_y5),
    .I0(1'b0),
    .I1(x17_y6),
    .I2(x16_y3),
    .I3(x17_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111100000101)
) lut_20_5 (
    .O(x20_y5),
    .I0(x17_y9),
    .I1(x18_y0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010001100000)
) lut_21_5 (
    .O(x21_y5),
    .I0(x18_y2),
    .I1(x19_y4),
    .I2(x18_y2),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010001001101)
) lut_22_5 (
    .O(x22_y5),
    .I0(x19_y5),
    .I1(x19_y10),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010001111110)
) lut_23_5 (
    .O(x23_y5),
    .I0(x21_y7),
    .I1(x21_y0),
    .I2(1'b0),
    .I3(x20_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010110110010)
) lut_24_5 (
    .O(x24_y5),
    .I0(x21_y0),
    .I1(x22_y0),
    .I2(x21_y0),
    .I3(x21_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001010010111)
) lut_25_5 (
    .O(x25_y5),
    .I0(x22_y9),
    .I1(x23_y8),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000011111011)
) lut_26_5 (
    .O(x26_y5),
    .I0(x24_y2),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x23_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000011100101)
) lut_27_5 (
    .O(x27_y5),
    .I0(x25_y3),
    .I1(x25_y8),
    .I2(1'b0),
    .I3(x25_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100011010001)
) lut_28_5 (
    .O(x28_y5),
    .I0(x25_y4),
    .I1(x25_y9),
    .I2(x25_y6),
    .I3(x25_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101000110101)
) lut_29_5 (
    .O(x29_y5),
    .I0(1'b0),
    .I1(x26_y0),
    .I2(x26_y10),
    .I3(x27_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100010110101)
) lut_30_5 (
    .O(x30_y5),
    .I0(x27_y7),
    .I1(x27_y8),
    .I2(x27_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100100011110)
) lut_31_5 (
    .O(x31_y5),
    .I0(1'b0),
    .I1(x29_y5),
    .I2(x29_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101000100110)
) lut_32_5 (
    .O(x32_y5),
    .I0(x29_y6),
    .I1(1'b0),
    .I2(x29_y5),
    .I3(x29_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101101100100)
) lut_33_5 (
    .O(x33_y5),
    .I0(1'b0),
    .I1(x30_y2),
    .I2(x31_y2),
    .I3(x31_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011111011110)
) lut_34_5 (
    .O(x34_y5),
    .I0(1'b0),
    .I1(x32_y1),
    .I2(x32_y7),
    .I3(x32_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011111111010)
) lut_35_5 (
    .O(x35_y5),
    .I0(x32_y6),
    .I1(x32_y7),
    .I2(x33_y8),
    .I3(x32_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101100010100)
) lut_36_5 (
    .O(x36_y5),
    .I0(x34_y4),
    .I1(1'b0),
    .I2(x34_y8),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010011111111)
) lut_37_5 (
    .O(x37_y5),
    .I0(x34_y10),
    .I1(x34_y5),
    .I2(x34_y10),
    .I3(x35_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001011000111)
) lut_38_5 (
    .O(x38_y5),
    .I0(1'b0),
    .I1(x35_y9),
    .I2(x36_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111001011011)
) lut_39_5 (
    .O(x39_y5),
    .I0(x37_y10),
    .I1(x37_y4),
    .I2(x36_y7),
    .I3(x36_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001000010010)
) lut_40_5 (
    .O(x40_y5),
    .I0(1'b0),
    .I1(x37_y8),
    .I2(x37_y8),
    .I3(x37_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110100010100)
) lut_41_5 (
    .O(x41_y5),
    .I0(x39_y4),
    .I1(x38_y4),
    .I2(x38_y6),
    .I3(x38_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001111001001)
) lut_42_5 (
    .O(x42_y5),
    .I0(x40_y3),
    .I1(x39_y2),
    .I2(x39_y3),
    .I3(x40_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111011110101)
) lut_43_5 (
    .O(x43_y5),
    .I0(x40_y10),
    .I1(x41_y0),
    .I2(x40_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011101111001)
) lut_44_5 (
    .O(x44_y5),
    .I0(x41_y3),
    .I1(x42_y1),
    .I2(1'b0),
    .I3(x41_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001111110001)
) lut_45_5 (
    .O(x45_y5),
    .I0(x43_y2),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x43_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101111111000)
) lut_46_5 (
    .O(x46_y5),
    .I0(1'b0),
    .I1(x44_y5),
    .I2(1'b0),
    .I3(x43_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010110010110)
) lut_47_5 (
    .O(x47_y5),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x44_y3),
    .I3(x44_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101100110111)
) lut_48_5 (
    .O(x48_y5),
    .I0(x46_y3),
    .I1(x45_y7),
    .I2(1'b0),
    .I3(x46_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001011110101)
) lut_49_5 (
    .O(x49_y5),
    .I0(1'b0),
    .I1(x47_y6),
    .I2(x46_y4),
    .I3(x46_y0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110011010101)
) lut_50_5 (
    .O(x50_y5),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x48_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010100100111)
) lut_51_5 (
    .O(x51_y5),
    .I0(x48_y4),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110011110011)
) lut_52_5 (
    .O(x52_y5),
    .I0(x50_y7),
    .I1(x49_y5),
    .I2(x49_y6),
    .I3(x50_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010000100000)
) lut_53_5 (
    .O(x53_y5),
    .I0(x51_y8),
    .I1(x51_y5),
    .I2(1'b0),
    .I3(x50_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010111010011)
) lut_54_5 (
    .O(x54_y5),
    .I0(1'b0),
    .I1(x52_y3),
    .I2(x51_y0),
    .I3(x52_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101111000110)
) lut_55_5 (
    .O(x55_y5),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x53_y8),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010100000000)
) lut_56_5 (
    .O(x56_y5),
    .I0(x53_y6),
    .I1(1'b0),
    .I2(x54_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011100001100)
) lut_57_5 (
    .O(x57_y5),
    .I0(x54_y1),
    .I1(x54_y5),
    .I2(x54_y2),
    .I3(x54_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110101100010)
) lut_58_5 (
    .O(x58_y5),
    .I0(x56_y0),
    .I1(x55_y7),
    .I2(x55_y7),
    .I3(x56_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011110100100)
) lut_59_5 (
    .O(x59_y5),
    .I0(x57_y1),
    .I1(1'b0),
    .I2(x57_y9),
    .I3(x57_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111010000011)
) lut_60_5 (
    .O(x60_y5),
    .I0(1'b0),
    .I1(x57_y10),
    .I2(1'b0),
    .I3(x58_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101111000110)
) lut_61_5 (
    .O(x61_y5),
    .I0(x59_y1),
    .I1(x59_y5),
    .I2(x59_y5),
    .I3(x59_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101111111110)
) lut_62_5 (
    .O(x62_y5),
    .I0(x60_y3),
    .I1(x59_y2),
    .I2(x60_y4),
    .I3(x59_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000111011111)
) lut_0_6 (
    .O(x0_y6),
    .I0(1'b0),
    .I1(in2),
    .I2(in6),
    .I3(in5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010001110100)
) lut_1_6 (
    .O(x1_y6),
    .I0(in3),
    .I1(in0),
    .I2(1'b0),
    .I3(in3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001001100111)
) lut_2_6 (
    .O(x2_y6),
    .I0(1'b0),
    .I1(in1),
    .I2(in5),
    .I3(in5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001110100111)
) lut_3_6 (
    .O(x3_y6),
    .I0(in2),
    .I1(in5),
    .I2(in4),
    .I3(x1_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100001101000)
) lut_4_6 (
    .O(x4_y6),
    .I0(x1_y9),
    .I1(x1_y2),
    .I2(x1_y8),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011110111001)
) lut_5_6 (
    .O(x5_y6),
    .I0(x2_y5),
    .I1(x3_y2),
    .I2(x2_y11),
    .I3(x2_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101110100011)
) lut_6_6 (
    .O(x6_y6),
    .I0(1'b0),
    .I1(x3_y3),
    .I2(x3_y7),
    .I3(x4_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000100001111)
) lut_7_6 (
    .O(x7_y6),
    .I0(x4_y4),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010001001110)
) lut_8_6 (
    .O(x8_y6),
    .I0(1'b0),
    .I1(x5_y7),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100111101000)
) lut_9_6 (
    .O(x9_y6),
    .I0(1'b0),
    .I1(x6_y8),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001010111011)
) lut_10_6 (
    .O(x10_y6),
    .I0(x8_y3),
    .I1(1'b0),
    .I2(x7_y3),
    .I3(x7_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011001110100)
) lut_11_6 (
    .O(x11_y6),
    .I0(1'b0),
    .I1(x8_y9),
    .I2(x9_y9),
    .I3(x8_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111010111110)
) lut_12_6 (
    .O(x12_y6),
    .I0(x10_y10),
    .I1(x10_y2),
    .I2(1'b0),
    .I3(x10_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101001100100)
) lut_13_6 (
    .O(x13_y6),
    .I0(1'b0),
    .I1(x10_y4),
    .I2(x11_y10),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001000110000)
) lut_14_6 (
    .O(x14_y6),
    .I0(x11_y2),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000100100100)
) lut_15_6 (
    .O(x15_y6),
    .I0(x12_y9),
    .I1(1'b0),
    .I2(x13_y1),
    .I3(x12_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000011011001)
) lut_16_6 (
    .O(x16_y6),
    .I0(x14_y5),
    .I1(x13_y11),
    .I2(x14_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000001111011)
) lut_17_6 (
    .O(x17_y6),
    .I0(1'b0),
    .I1(x15_y2),
    .I2(x15_y10),
    .I3(x15_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101010000101)
) lut_18_6 (
    .O(x18_y6),
    .I0(x16_y2),
    .I1(1'b0),
    .I2(x15_y8),
    .I3(x15_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111000110010)
) lut_19_6 (
    .O(x19_y6),
    .I0(x16_y4),
    .I1(x17_y6),
    .I2(1'b0),
    .I3(x16_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010010101100)
) lut_20_6 (
    .O(x20_y6),
    .I0(x17_y2),
    .I1(x18_y4),
    .I2(x17_y7),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101101101011)
) lut_21_6 (
    .O(x21_y6),
    .I0(x18_y3),
    .I1(x18_y3),
    .I2(x19_y4),
    .I3(x19_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000011011110)
) lut_22_6 (
    .O(x22_y6),
    .I0(x20_y6),
    .I1(x20_y3),
    .I2(x20_y7),
    .I3(x19_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011111111000)
) lut_23_6 (
    .O(x23_y6),
    .I0(x20_y9),
    .I1(x20_y3),
    .I2(x20_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100010111001)
) lut_24_6 (
    .O(x24_y6),
    .I0(x22_y5),
    .I1(x22_y6),
    .I2(1'b0),
    .I3(x21_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101101000011)
) lut_25_6 (
    .O(x25_y6),
    .I0(x22_y4),
    .I1(x22_y5),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000101100000)
) lut_26_6 (
    .O(x26_y6),
    .I0(x24_y3),
    .I1(x23_y7),
    .I2(x23_y1),
    .I3(x24_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011100101000)
) lut_27_6 (
    .O(x27_y6),
    .I0(x24_y7),
    .I1(1'b0),
    .I2(x25_y3),
    .I3(x25_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011010111011)
) lut_28_6 (
    .O(x28_y6),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x25_y1),
    .I3(x25_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111011000100)
) lut_29_6 (
    .O(x29_y6),
    .I0(x26_y5),
    .I1(x27_y7),
    .I2(1'b0),
    .I3(x26_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010011110011)
) lut_30_6 (
    .O(x30_y6),
    .I0(x27_y7),
    .I1(x28_y2),
    .I2(x28_y11),
    .I3(x28_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111100010001)
) lut_31_6 (
    .O(x31_y6),
    .I0(x29_y5),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100101000111)
) lut_32_6 (
    .O(x32_y6),
    .I0(x30_y4),
    .I1(1'b0),
    .I2(x30_y11),
    .I3(x29_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011011101000)
) lut_33_6 (
    .O(x33_y6),
    .I0(x31_y7),
    .I1(1'b0),
    .I2(x31_y1),
    .I3(x31_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001111111111)
) lut_34_6 (
    .O(x34_y6),
    .I0(x32_y5),
    .I1(1'b0),
    .I2(x32_y1),
    .I3(x32_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010001110010)
) lut_35_6 (
    .O(x35_y6),
    .I0(x32_y4),
    .I1(x33_y7),
    .I2(x33_y1),
    .I3(x32_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010111101101)
) lut_36_6 (
    .O(x36_y6),
    .I0(x34_y4),
    .I1(x33_y1),
    .I2(x33_y7),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011110101110)
) lut_37_6 (
    .O(x37_y6),
    .I0(x34_y6),
    .I1(1'b0),
    .I2(x35_y2),
    .I3(x35_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110101100011)
) lut_38_6 (
    .O(x38_y6),
    .I0(x35_y5),
    .I1(1'b0),
    .I2(x35_y7),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011111101010)
) lut_39_6 (
    .O(x39_y6),
    .I0(x37_y9),
    .I1(x36_y5),
    .I2(x37_y9),
    .I3(x36_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110001111010)
) lut_40_6 (
    .O(x40_y6),
    .I0(x38_y9),
    .I1(x37_y2),
    .I2(x38_y4),
    .I3(x38_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101010100011)
) lut_41_6 (
    .O(x41_y6),
    .I0(x39_y2),
    .I1(x38_y9),
    .I2(x38_y3),
    .I3(x38_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010110100101)
) lut_42_6 (
    .O(x42_y6),
    .I0(x40_y5),
    .I1(x39_y1),
    .I2(x40_y5),
    .I3(x39_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110111011111)
) lut_43_6 (
    .O(x43_y6),
    .I0(1'b0),
    .I1(x41_y10),
    .I2(x40_y1),
    .I3(x40_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101110100110)
) lut_44_6 (
    .O(x44_y6),
    .I0(x41_y10),
    .I1(1'b0),
    .I2(x41_y7),
    .I3(x41_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010010110111)
) lut_45_6 (
    .O(x45_y6),
    .I0(x42_y5),
    .I1(x43_y2),
    .I2(1'b0),
    .I3(x42_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110001101011)
) lut_46_6 (
    .O(x46_y6),
    .I0(1'b0),
    .I1(x43_y8),
    .I2(x44_y11),
    .I3(x43_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100010011100)
) lut_47_6 (
    .O(x47_y6),
    .I0(1'b0),
    .I1(x45_y4),
    .I2(x45_y8),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111111000001)
) lut_48_6 (
    .O(x48_y6),
    .I0(x45_y7),
    .I1(x45_y2),
    .I2(x46_y3),
    .I3(x46_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000101010000)
) lut_49_6 (
    .O(x49_y6),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x47_y9),
    .I3(x46_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110110010101)
) lut_50_6 (
    .O(x50_y6),
    .I0(1'b0),
    .I1(x47_y6),
    .I2(x47_y8),
    .I3(x48_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010000010000)
) lut_51_6 (
    .O(x51_y6),
    .I0(x48_y10),
    .I1(x49_y5),
    .I2(x49_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101100001001)
) lut_52_6 (
    .O(x52_y6),
    .I0(x49_y6),
    .I1(x50_y1),
    .I2(x49_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000101010010)
) lut_53_6 (
    .O(x53_y6),
    .I0(1'b0),
    .I1(x51_y3),
    .I2(x51_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100111110100)
) lut_54_6 (
    .O(x54_y6),
    .I0(x51_y5),
    .I1(x52_y6),
    .I2(1'b0),
    .I3(x51_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101010101011)
) lut_55_6 (
    .O(x55_y6),
    .I0(x52_y4),
    .I1(x52_y4),
    .I2(x52_y9),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001011000010)
) lut_56_6 (
    .O(x56_y6),
    .I0(1'b0),
    .I1(x53_y2),
    .I2(x54_y1),
    .I3(x53_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111011000101)
) lut_57_6 (
    .O(x57_y6),
    .I0(x54_y1),
    .I1(x55_y4),
    .I2(1'b0),
    .I3(x55_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110011110100)
) lut_58_6 (
    .O(x58_y6),
    .I0(x56_y3),
    .I1(x55_y6),
    .I2(x56_y11),
    .I3(x55_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001101000110)
) lut_59_6 (
    .O(x59_y6),
    .I0(x57_y9),
    .I1(1'b0),
    .I2(x57_y1),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000110110111)
) lut_60_6 (
    .O(x60_y6),
    .I0(x57_y4),
    .I1(1'b0),
    .I2(x58_y8),
    .I3(x57_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010100111100)
) lut_61_6 (
    .O(x61_y6),
    .I0(x59_y7),
    .I1(x59_y11),
    .I2(x58_y9),
    .I3(x59_y1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110001101001)
) lut_62_6 (
    .O(x62_y6),
    .I0(x60_y7),
    .I1(1'b0),
    .I2(x59_y1),
    .I3(x59_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001001011101)
) lut_0_7 (
    .O(x0_y7),
    .I0(in5),
    .I1(in5),
    .I2(in1),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111101101111)
) lut_1_7 (
    .O(x1_y7),
    .I0(in5),
    .I1(in4),
    .I2(in1),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001100110010)
) lut_2_7 (
    .O(x2_y7),
    .I0(in6),
    .I1(in7),
    .I2(in2),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010100111111)
) lut_3_7 (
    .O(x3_y7),
    .I0(in1),
    .I1(in5),
    .I2(in3),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101010110000)
) lut_4_7 (
    .O(x4_y7),
    .I0(x2_y6),
    .I1(x2_y11),
    .I2(1'b0),
    .I3(x1_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111100011111)
) lut_5_7 (
    .O(x5_y7),
    .I0(x2_y3),
    .I1(1'b0),
    .I2(x3_y8),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001110001101)
) lut_6_7 (
    .O(x6_y7),
    .I0(x4_y12),
    .I1(x4_y7),
    .I2(x4_y6),
    .I3(x4_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100100010011)
) lut_7_7 (
    .O(x7_y7),
    .I0(1'b0),
    .I1(x4_y6),
    .I2(x5_y3),
    .I3(x5_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100010001011)
) lut_8_7 (
    .O(x8_y7),
    .I0(x6_y6),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x6_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110111010110)
) lut_9_7 (
    .O(x9_y7),
    .I0(x7_y10),
    .I1(x6_y4),
    .I2(1'b0),
    .I3(x6_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000101000110)
) lut_10_7 (
    .O(x10_y7),
    .I0(1'b0),
    .I1(x7_y12),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110110111001)
) lut_11_7 (
    .O(x11_y7),
    .I0(x8_y7),
    .I1(x8_y7),
    .I2(1'b0),
    .I3(x8_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101010010111)
) lut_12_7 (
    .O(x12_y7),
    .I0(x9_y5),
    .I1(x9_y4),
    .I2(x10_y8),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010101111101)
) lut_13_7 (
    .O(x13_y7),
    .I0(x11_y10),
    .I1(x11_y3),
    .I2(x11_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111010101010)
) lut_14_7 (
    .O(x14_y7),
    .I0(x12_y6),
    .I1(x12_y10),
    .I2(x11_y7),
    .I3(x11_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011110001000)
) lut_15_7 (
    .O(x15_y7),
    .I0(x12_y10),
    .I1(1'b0),
    .I2(x13_y11),
    .I3(x13_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111001000110)
) lut_16_7 (
    .O(x16_y7),
    .I0(x14_y11),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x13_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001010001011)
) lut_17_7 (
    .O(x17_y7),
    .I0(x15_y8),
    .I1(x14_y2),
    .I2(x15_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100010001000)
) lut_18_7 (
    .O(x18_y7),
    .I0(x16_y3),
    .I1(x16_y7),
    .I2(x15_y12),
    .I3(x15_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010100001010)
) lut_19_7 (
    .O(x19_y7),
    .I0(x16_y9),
    .I1(x17_y11),
    .I2(x17_y5),
    .I3(x16_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000011001011)
) lut_20_7 (
    .O(x20_y7),
    .I0(x17_y12),
    .I1(x17_y7),
    .I2(x18_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111100111001)
) lut_21_7 (
    .O(x21_y7),
    .I0(x18_y6),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x18_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101100010001)
) lut_22_7 (
    .O(x22_y7),
    .I0(x19_y11),
    .I1(x20_y8),
    .I2(x19_y11),
    .I3(x20_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100010010101)
) lut_23_7 (
    .O(x23_y7),
    .I0(1'b0),
    .I1(x20_y6),
    .I2(x21_y12),
    .I3(x21_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100001001100)
) lut_24_7 (
    .O(x24_y7),
    .I0(x22_y3),
    .I1(x22_y7),
    .I2(x22_y6),
    .I3(x21_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101101111010)
) lut_25_7 (
    .O(x25_y7),
    .I0(x22_y4),
    .I1(1'b0),
    .I2(x22_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011100111011)
) lut_26_7 (
    .O(x26_y7),
    .I0(x24_y6),
    .I1(x23_y11),
    .I2(x24_y10),
    .I3(x24_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101111010110)
) lut_27_7 (
    .O(x27_y7),
    .I0(x24_y9),
    .I1(x25_y4),
    .I2(x24_y8),
    .I3(x25_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111111100011)
) lut_28_7 (
    .O(x28_y7),
    .I0(x26_y6),
    .I1(x25_y5),
    .I2(x25_y12),
    .I3(x26_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011011110110)
) lut_29_7 (
    .O(x29_y7),
    .I0(x27_y6),
    .I1(x26_y11),
    .I2(x27_y2),
    .I3(x27_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000101000011)
) lut_30_7 (
    .O(x30_y7),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x27_y3),
    .I3(x28_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100001101010)
) lut_31_7 (
    .O(x31_y7),
    .I0(1'b0),
    .I1(x28_y12),
    .I2(x29_y12),
    .I3(x29_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101000010010)
) lut_32_7 (
    .O(x32_y7),
    .I0(x30_y2),
    .I1(1'b0),
    .I2(x30_y6),
    .I3(x30_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110110110011)
) lut_33_7 (
    .O(x33_y7),
    .I0(x31_y8),
    .I1(x30_y2),
    .I2(x31_y6),
    .I3(x30_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011100011000)
) lut_34_7 (
    .O(x34_y7),
    .I0(x31_y12),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x32_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011010111000)
) lut_35_7 (
    .O(x35_y7),
    .I0(x32_y12),
    .I1(x32_y4),
    .I2(x32_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001101010001)
) lut_36_7 (
    .O(x36_y7),
    .I0(x33_y11),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x34_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001110100100)
) lut_37_7 (
    .O(x37_y7),
    .I0(x34_y2),
    .I1(x35_y5),
    .I2(1'b0),
    .I3(x35_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011100100111)
) lut_38_7 (
    .O(x38_y7),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x35_y12),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010100010111)
) lut_39_7 (
    .O(x39_y7),
    .I0(x36_y10),
    .I1(x37_y10),
    .I2(x37_y4),
    .I3(x36_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110100011010)
) lut_40_7 (
    .O(x40_y7),
    .I0(x37_y12),
    .I1(x38_y6),
    .I2(x38_y7),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110001000001)
) lut_41_7 (
    .O(x41_y7),
    .I0(x38_y5),
    .I1(x38_y9),
    .I2(x39_y6),
    .I3(x38_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000110001110)
) lut_42_7 (
    .O(x42_y7),
    .I0(1'b0),
    .I1(x39_y2),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011110000111)
) lut_43_7 (
    .O(x43_y7),
    .I0(1'b0),
    .I1(x41_y2),
    .I2(x41_y4),
    .I3(x41_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000111000010)
) lut_44_7 (
    .O(x44_y7),
    .I0(x42_y6),
    .I1(x41_y3),
    .I2(1'b0),
    .I3(x41_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111110111001)
) lut_45_7 (
    .O(x45_y7),
    .I0(x43_y4),
    .I1(x43_y4),
    .I2(x42_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100100000001)
) lut_46_7 (
    .O(x46_y7),
    .I0(x43_y9),
    .I1(x44_y2),
    .I2(x43_y12),
    .I3(x43_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100001000011)
) lut_47_7 (
    .O(x47_y7),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x44_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000110101110)
) lut_48_7 (
    .O(x48_y7),
    .I0(x45_y5),
    .I1(x46_y7),
    .I2(x46_y7),
    .I3(x45_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100011110111)
) lut_49_7 (
    .O(x49_y7),
    .I0(x46_y3),
    .I1(1'b0),
    .I2(x46_y7),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001011100011)
) lut_50_7 (
    .O(x50_y7),
    .I0(x48_y4),
    .I1(x47_y5),
    .I2(x47_y5),
    .I3(x48_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110110001100)
) lut_51_7 (
    .O(x51_y7),
    .I0(1'b0),
    .I1(x48_y12),
    .I2(x49_y9),
    .I3(x48_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000010111101)
) lut_52_7 (
    .O(x52_y7),
    .I0(x49_y3),
    .I1(x50_y12),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010110011001)
) lut_53_7 (
    .O(x53_y7),
    .I0(x51_y6),
    .I1(1'b0),
    .I2(x51_y8),
    .I3(x51_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111011001111)
) lut_54_7 (
    .O(x54_y7),
    .I0(x51_y8),
    .I1(x51_y5),
    .I2(x52_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110011101111)
) lut_55_7 (
    .O(x55_y7),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x53_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101001001101)
) lut_56_7 (
    .O(x56_y7),
    .I0(1'b0),
    .I1(x54_y3),
    .I2(x53_y11),
    .I3(x54_y3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000100101100)
) lut_57_7 (
    .O(x57_y7),
    .I0(x54_y10),
    .I1(x55_y7),
    .I2(x55_y7),
    .I3(x55_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010100100011)
) lut_58_7 (
    .O(x58_y7),
    .I0(x56_y3),
    .I1(1'b0),
    .I2(x55_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101011100101)
) lut_59_7 (
    .O(x59_y7),
    .I0(1'b0),
    .I1(x57_y4),
    .I2(x57_y5),
    .I3(x56_y2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011110010110)
) lut_60_7 (
    .O(x60_y7),
    .I0(x58_y12),
    .I1(x57_y8),
    .I2(x57_y10),
    .I3(x58_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111101011011)
) lut_61_7 (
    .O(x61_y7),
    .I0(x59_y11),
    .I1(x58_y2),
    .I2(1'b0),
    .I3(x58_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100111101100)
) lut_62_7 (
    .O(x62_y7),
    .I0(1'b0),
    .I1(x60_y12),
    .I2(x60_y12),
    .I3(x59_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110100011110)
) lut_0_8 (
    .O(x0_y8),
    .I0(in8),
    .I1(in6),
    .I2(in1),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011111000010)
) lut_1_8 (
    .O(x1_y8),
    .I0(in4),
    .I1(in8),
    .I2(in1),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011100101101)
) lut_2_8 (
    .O(x2_y8),
    .I0(1'b0),
    .I1(in5),
    .I2(in7),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100000000001)
) lut_3_8 (
    .O(x3_y8),
    .I0(in3),
    .I1(in2),
    .I2(in7),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001011011100)
) lut_4_8 (
    .O(x4_y8),
    .I0(x1_y12),
    .I1(x1_y3),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001110011010)
) lut_5_8 (
    .O(x5_y8),
    .I0(1'b0),
    .I1(x3_y12),
    .I2(x3_y7),
    .I3(x3_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100111001110)
) lut_6_8 (
    .O(x6_y8),
    .I0(x4_y12),
    .I1(x4_y6),
    .I2(x3_y10),
    .I3(x4_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101101011110)
) lut_7_8 (
    .O(x7_y8),
    .I0(x5_y11),
    .I1(x4_y7),
    .I2(x5_y9),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101000001000)
) lut_8_8 (
    .O(x8_y8),
    .I0(x5_y5),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101001111101)
) lut_9_8 (
    .O(x9_y8),
    .I0(x7_y12),
    .I1(x6_y12),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000111001111)
) lut_10_8 (
    .O(x10_y8),
    .I0(x7_y5),
    .I1(x7_y5),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001100101101)
) lut_11_8 (
    .O(x11_y8),
    .I0(x9_y7),
    .I1(x9_y6),
    .I2(x9_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101111100100)
) lut_12_8 (
    .O(x12_y8),
    .I0(1'b0),
    .I1(x10_y7),
    .I2(x9_y4),
    .I3(x10_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010011100101)
) lut_13_8 (
    .O(x13_y8),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x10_y11),
    .I3(x11_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010010101100)
) lut_14_8 (
    .O(x14_y8),
    .I0(x11_y5),
    .I1(x11_y3),
    .I2(x11_y13),
    .I3(x12_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010001111000)
) lut_15_8 (
    .O(x15_y8),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x13_y11),
    .I3(x12_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000010010110)
) lut_16_8 (
    .O(x16_y8),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x13_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010000011100)
) lut_17_8 (
    .O(x17_y8),
    .I0(x15_y9),
    .I1(x14_y11),
    .I2(x14_y7),
    .I3(x14_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010100011111)
) lut_18_8 (
    .O(x18_y8),
    .I0(1'b0),
    .I1(x16_y8),
    .I2(x15_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000001011111)
) lut_19_8 (
    .O(x19_y8),
    .I0(x16_y3),
    .I1(x16_y3),
    .I2(x17_y5),
    .I3(x16_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110011110110)
) lut_20_8 (
    .O(x20_y8),
    .I0(x18_y8),
    .I1(x18_y5),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101110000001)
) lut_21_8 (
    .O(x21_y8),
    .I0(x19_y9),
    .I1(x19_y4),
    .I2(x19_y8),
    .I3(x18_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111010111100)
) lut_22_8 (
    .O(x22_y8),
    .I0(x20_y10),
    .I1(x20_y13),
    .I2(x20_y5),
    .I3(x19_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111111011000)
) lut_23_8 (
    .O(x23_y8),
    .I0(x21_y3),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010011110000)
) lut_24_8 (
    .O(x24_y8),
    .I0(1'b0),
    .I1(x21_y6),
    .I2(x22_y8),
    .I3(x21_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010010001011)
) lut_25_8 (
    .O(x25_y8),
    .I0(x23_y7),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x22_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001000110110)
) lut_26_8 (
    .O(x26_y8),
    .I0(x23_y12),
    .I1(1'b0),
    .I2(x24_y5),
    .I3(x24_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010000011011)
) lut_27_8 (
    .O(x27_y8),
    .I0(x24_y13),
    .I1(1'b0),
    .I2(x24_y3),
    .I3(x24_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100100101011)
) lut_28_8 (
    .O(x28_y8),
    .I0(1'b0),
    .I1(x26_y4),
    .I2(x25_y10),
    .I3(x25_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010011000011)
) lut_29_8 (
    .O(x29_y8),
    .I0(1'b0),
    .I1(x27_y5),
    .I2(x27_y11),
    .I3(x26_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001101100000)
) lut_30_8 (
    .O(x30_y8),
    .I0(x28_y12),
    .I1(x27_y6),
    .I2(x28_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101100001101)
) lut_31_8 (
    .O(x31_y8),
    .I0(x29_y9),
    .I1(1'b0),
    .I2(x29_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111011100110)
) lut_32_8 (
    .O(x32_y8),
    .I0(x30_y3),
    .I1(x30_y6),
    .I2(1'b0),
    .I3(x30_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100111010011)
) lut_33_8 (
    .O(x33_y8),
    .I0(x30_y8),
    .I1(1'b0),
    .I2(x30_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001011100011)
) lut_34_8 (
    .O(x34_y8),
    .I0(x32_y9),
    .I1(x32_y10),
    .I2(x32_y5),
    .I3(x31_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011011101111)
) lut_35_8 (
    .O(x35_y8),
    .I0(1'b0),
    .I1(x32_y12),
    .I2(x33_y11),
    .I3(x32_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010100011111)
) lut_36_8 (
    .O(x36_y8),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x34_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000100010110)
) lut_37_8 (
    .O(x37_y8),
    .I0(x34_y3),
    .I1(x35_y6),
    .I2(x34_y10),
    .I3(x34_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111111110100)
) lut_38_8 (
    .O(x38_y8),
    .I0(x35_y6),
    .I1(x35_y8),
    .I2(1'b0),
    .I3(x36_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000110101011)
) lut_39_8 (
    .O(x39_y8),
    .I0(1'b0),
    .I1(x37_y4),
    .I2(x37_y6),
    .I3(x36_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001111100010)
) lut_40_8 (
    .O(x40_y8),
    .I0(x38_y3),
    .I1(x37_y11),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011110001101)
) lut_41_8 (
    .O(x41_y8),
    .I0(x39_y12),
    .I1(x38_y7),
    .I2(1'b0),
    .I3(x38_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001100010101)
) lut_42_8 (
    .O(x42_y8),
    .I0(x40_y12),
    .I1(x40_y12),
    .I2(1'b0),
    .I3(x40_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110110111000)
) lut_43_8 (
    .O(x43_y8),
    .I0(x41_y6),
    .I1(x40_y8),
    .I2(1'b0),
    .I3(x40_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100101010100)
) lut_44_8 (
    .O(x44_y8),
    .I0(x42_y9),
    .I1(x42_y12),
    .I2(x42_y4),
    .I3(x42_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010011001010)
) lut_45_8 (
    .O(x45_y8),
    .I0(x42_y7),
    .I1(x42_y6),
    .I2(1'b0),
    .I3(x43_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000001000000)
) lut_46_8 (
    .O(x46_y8),
    .I0(x44_y11),
    .I1(1'b0),
    .I2(x43_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011010111110)
) lut_47_8 (
    .O(x47_y8),
    .I0(x44_y8),
    .I1(1'b0),
    .I2(x44_y4),
    .I3(x44_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010010101000)
) lut_48_8 (
    .O(x48_y8),
    .I0(x45_y3),
    .I1(x46_y3),
    .I2(x46_y3),
    .I3(x45_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101011110110)
) lut_49_8 (
    .O(x49_y8),
    .I0(1'b0),
    .I1(x47_y10),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101011111000)
) lut_50_8 (
    .O(x50_y8),
    .I0(x48_y9),
    .I1(x47_y12),
    .I2(1'b0),
    .I3(x47_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000111101110)
) lut_51_8 (
    .O(x51_y8),
    .I0(x49_y7),
    .I1(x49_y11),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000000001111)
) lut_52_8 (
    .O(x52_y8),
    .I0(x50_y4),
    .I1(1'b0),
    .I2(x50_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111010010110)
) lut_53_8 (
    .O(x53_y8),
    .I0(x51_y5),
    .I1(x51_y5),
    .I2(1'b0),
    .I3(x50_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000000101110)
) lut_54_8 (
    .O(x54_y8),
    .I0(1'b0),
    .I1(x52_y9),
    .I2(x51_y9),
    .I3(x51_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001101100000)
) lut_55_8 (
    .O(x55_y8),
    .I0(x53_y6),
    .I1(x52_y6),
    .I2(1'b0),
    .I3(x53_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000100101000)
) lut_56_8 (
    .O(x56_y8),
    .I0(x54_y13),
    .I1(x54_y7),
    .I2(x54_y3),
    .I3(x53_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010101010001)
) lut_57_8 (
    .O(x57_y8),
    .I0(x54_y7),
    .I1(x55_y7),
    .I2(x54_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110111111100)
) lut_58_8 (
    .O(x58_y8),
    .I0(1'b0),
    .I1(x55_y9),
    .I2(x56_y11),
    .I3(x55_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101011101110)
) lut_59_8 (
    .O(x59_y8),
    .I0(x57_y13),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x56_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101010011010)
) lut_60_8 (
    .O(x60_y8),
    .I0(1'b0),
    .I1(x57_y13),
    .I2(x58_y13),
    .I3(x58_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111101110111)
) lut_61_8 (
    .O(x61_y8),
    .I0(x59_y11),
    .I1(x59_y3),
    .I2(x58_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010011100010)
) lut_62_8 (
    .O(x62_y8),
    .I0(x60_y5),
    .I1(1'b0),
    .I2(x59_y6),
    .I3(x60_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110110100101)
) lut_0_9 (
    .O(x0_y9),
    .I0(in7),
    .I1(in7),
    .I2(in6),
    .I3(in4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101100010000)
) lut_1_9 (
    .O(x1_y9),
    .I0(in2),
    .I1(in4),
    .I2(in5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000001101011)
) lut_2_9 (
    .O(x2_y9),
    .I0(in9),
    .I1(in4),
    .I2(in6),
    .I3(in7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100101011100)
) lut_3_9 (
    .O(x3_y9),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100011110011)
) lut_4_9 (
    .O(x4_y9),
    .I0(x2_y5),
    .I1(x2_y4),
    .I2(x1_y9),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111011001110)
) lut_5_9 (
    .O(x5_y9),
    .I0(1'b0),
    .I1(x2_y5),
    .I2(x3_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010111111101)
) lut_6_9 (
    .O(x6_y9),
    .I0(x3_y13),
    .I1(x4_y12),
    .I2(x3_y8),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011010110111)
) lut_7_9 (
    .O(x7_y9),
    .I0(x5_y6),
    .I1(x5_y10),
    .I2(x4_y9),
    .I3(x4_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011000010101)
) lut_8_9 (
    .O(x8_y9),
    .I0(x5_y7),
    .I1(x5_y6),
    .I2(x5_y7),
    .I3(x5_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110001001101)
) lut_9_9 (
    .O(x9_y9),
    .I0(x6_y7),
    .I1(1'b0),
    .I2(x5_y7),
    .I3(x5_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010001101100)
) lut_10_9 (
    .O(x10_y9),
    .I0(1'b0),
    .I1(x7_y6),
    .I2(x8_y10),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110000100010)
) lut_11_9 (
    .O(x11_y9),
    .I0(x8_y8),
    .I1(x8_y4),
    .I2(x8_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110110110000)
) lut_12_9 (
    .O(x12_y9),
    .I0(x10_y9),
    .I1(x10_y12),
    .I2(1'b0),
    .I3(x9_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010010111111)
) lut_13_9 (
    .O(x13_y9),
    .I0(x11_y13),
    .I1(x11_y14),
    .I2(x11_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100001101101)
) lut_14_9 (
    .O(x14_y9),
    .I0(x11_y13),
    .I1(x12_y4),
    .I2(x11_y6),
    .I3(x11_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001000010010)
) lut_15_9 (
    .O(x15_y9),
    .I0(x12_y9),
    .I1(x12_y5),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000000001010)
) lut_16_9 (
    .O(x16_y9),
    .I0(x13_y6),
    .I1(x13_y6),
    .I2(x13_y6),
    .I3(x13_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000100100011)
) lut_17_9 (
    .O(x17_y9),
    .I0(x14_y5),
    .I1(x14_y13),
    .I2(x15_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010001001001)
) lut_18_9 (
    .O(x18_y9),
    .I0(x16_y10),
    .I1(x15_y13),
    .I2(x15_y5),
    .I3(x15_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110010000001)
) lut_19_9 (
    .O(x19_y9),
    .I0(1'b0),
    .I1(x16_y6),
    .I2(x16_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001111001011)
) lut_20_9 (
    .O(x20_y9),
    .I0(x17_y8),
    .I1(x18_y10),
    .I2(1'b0),
    .I3(x17_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010111101110)
) lut_21_9 (
    .O(x21_y9),
    .I0(x19_y11),
    .I1(1'b0),
    .I2(x18_y5),
    .I3(x19_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101010010101)
) lut_22_9 (
    .O(x22_y9),
    .I0(1'b0),
    .I1(x20_y7),
    .I2(x20_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001100100101)
) lut_23_9 (
    .O(x23_y9),
    .I0(x20_y4),
    .I1(x21_y6),
    .I2(x20_y7),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101111100010)
) lut_24_9 (
    .O(x24_y9),
    .I0(1'b0),
    .I1(x22_y9),
    .I2(x22_y5),
    .I3(x21_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101101010011)
) lut_25_9 (
    .O(x25_y9),
    .I0(1'b0),
    .I1(x22_y6),
    .I2(x23_y5),
    .I3(x22_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000001101100)
) lut_26_9 (
    .O(x26_y9),
    .I0(x24_y5),
    .I1(x23_y14),
    .I2(x23_y13),
    .I3(x24_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000110100100)
) lut_27_9 (
    .O(x27_y9),
    .I0(x25_y12),
    .I1(x25_y8),
    .I2(x25_y14),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011011111000)
) lut_28_9 (
    .O(x28_y9),
    .I0(x26_y12),
    .I1(x25_y9),
    .I2(x25_y9),
    .I3(x25_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000011011100)
) lut_29_9 (
    .O(x29_y9),
    .I0(x27_y7),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x26_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000101001011)
) lut_30_9 (
    .O(x30_y9),
    .I0(x28_y8),
    .I1(1'b0),
    .I2(x28_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100000101100)
) lut_31_9 (
    .O(x31_y9),
    .I0(x29_y13),
    .I1(x28_y9),
    .I2(x29_y12),
    .I3(x29_y4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111100101001)
) lut_32_9 (
    .O(x32_y9),
    .I0(x30_y4),
    .I1(x30_y13),
    .I2(1'b0),
    .I3(x29_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100110000001)
) lut_33_9 (
    .O(x33_y9),
    .I0(x31_y13),
    .I1(1'b0),
    .I2(x30_y10),
    .I3(x30_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100111000110)
) lut_34_9 (
    .O(x34_y9),
    .I0(x31_y11),
    .I1(x32_y14),
    .I2(x31_y5),
    .I3(x31_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111101000100)
) lut_35_9 (
    .O(x35_y9),
    .I0(x32_y10),
    .I1(x32_y7),
    .I2(x33_y6),
    .I3(x32_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101011100000)
) lut_36_9 (
    .O(x36_y9),
    .I0(x33_y10),
    .I1(x34_y11),
    .I2(x33_y9),
    .I3(x34_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011100011110)
) lut_37_9 (
    .O(x37_y9),
    .I0(1'b0),
    .I1(x34_y14),
    .I2(x34_y11),
    .I3(x34_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010010110110)
) lut_38_9 (
    .O(x38_y9),
    .I0(x36_y5),
    .I1(x35_y9),
    .I2(x35_y5),
    .I3(x35_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000010111110)
) lut_39_9 (
    .O(x39_y9),
    .I0(1'b0),
    .I1(x36_y13),
    .I2(x36_y11),
    .I3(x37_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011001010110)
) lut_40_9 (
    .O(x40_y9),
    .I0(x37_y14),
    .I1(1'b0),
    .I2(x38_y9),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111001001010)
) lut_41_9 (
    .O(x41_y9),
    .I0(x39_y5),
    .I1(1'b0),
    .I2(x39_y8),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001111001111)
) lut_42_9 (
    .O(x42_y9),
    .I0(x40_y6),
    .I1(x40_y5),
    .I2(x40_y7),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101110000100)
) lut_43_9 (
    .O(x43_y9),
    .I0(x40_y14),
    .I1(x41_y14),
    .I2(1'b0),
    .I3(x40_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101110110101)
) lut_44_9 (
    .O(x44_y9),
    .I0(x42_y4),
    .I1(x41_y14),
    .I2(1'b0),
    .I3(x42_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100111111110)
) lut_45_9 (
    .O(x45_y9),
    .I0(x42_y7),
    .I1(x42_y7),
    .I2(x43_y7),
    .I3(x42_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101000001101)
) lut_46_9 (
    .O(x46_y9),
    .I0(x43_y4),
    .I1(1'b0),
    .I2(x43_y13),
    .I3(x44_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011101101101)
) lut_47_9 (
    .O(x47_y9),
    .I0(x45_y6),
    .I1(x45_y9),
    .I2(x44_y5),
    .I3(x45_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101111111010)
) lut_48_9 (
    .O(x48_y9),
    .I0(x45_y13),
    .I1(x45_y5),
    .I2(x45_y6),
    .I3(x45_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101010000010)
) lut_49_9 (
    .O(x49_y9),
    .I0(x47_y13),
    .I1(x46_y8),
    .I2(1'b0),
    .I3(x46_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101100101011)
) lut_50_9 (
    .O(x50_y9),
    .I0(x48_y5),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110001011000)
) lut_51_9 (
    .O(x51_y9),
    .I0(x49_y9),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011010111111)
) lut_52_9 (
    .O(x52_y9),
    .I0(x50_y5),
    .I1(x49_y6),
    .I2(1'b0),
    .I3(x49_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010101001110)
) lut_53_9 (
    .O(x53_y9),
    .I0(1'b0),
    .I1(x51_y13),
    .I2(x50_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000110100101)
) lut_54_9 (
    .O(x54_y9),
    .I0(1'b0),
    .I1(x51_y5),
    .I2(x52_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110100000111)
) lut_55_9 (
    .O(x55_y9),
    .I0(x53_y12),
    .I1(x53_y6),
    .I2(x53_y10),
    .I3(x52_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111110001011)
) lut_56_9 (
    .O(x56_y9),
    .I0(x54_y8),
    .I1(x54_y11),
    .I2(x54_y12),
    .I3(x53_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111010101110)
) lut_57_9 (
    .O(x57_y9),
    .I0(1'b0),
    .I1(x55_y11),
    .I2(x55_y10),
    .I3(x55_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000011001000)
) lut_58_9 (
    .O(x58_y9),
    .I0(x55_y6),
    .I1(x56_y8),
    .I2(x55_y10),
    .I3(x56_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001101011001)
) lut_59_9 (
    .O(x59_y9),
    .I0(x57_y11),
    .I1(x57_y8),
    .I2(x57_y13),
    .I3(x56_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100101001001)
) lut_60_9 (
    .O(x60_y9),
    .I0(x58_y10),
    .I1(x58_y6),
    .I2(x58_y7),
    .I3(x58_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010101011011)
) lut_61_9 (
    .O(x61_y9),
    .I0(x58_y7),
    .I1(x59_y8),
    .I2(x58_y13),
    .I3(x58_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010110001010)
) lut_62_9 (
    .O(x62_y9),
    .I0(x59_y13),
    .I1(x60_y14),
    .I2(x59_y10),
    .I3(x60_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100011111000)
) lut_0_10 (
    .O(x0_y10),
    .I0(in9),
    .I1(in5),
    .I2(in5),
    .I3(in7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001011101011)
) lut_1_10 (
    .O(x1_y10),
    .I0(in1),
    .I1(1'b0),
    .I2(in5),
    .I3(in4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011011100100)
) lut_2_10 (
    .O(x2_y10),
    .I0(1'b0),
    .I1(in4),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001100000100)
) lut_3_10 (
    .O(x3_y10),
    .I0(in8),
    .I1(in3),
    .I2(in8),
    .I3(in5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010001111010)
) lut_4_10 (
    .O(x4_y10),
    .I0(x2_y7),
    .I1(x1_y12),
    .I2(x1_y9),
    .I3(x1_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110101011100)
) lut_5_10 (
    .O(x5_y10),
    .I0(x2_y15),
    .I1(x3_y15),
    .I2(x3_y6),
    .I3(x2_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001000111100)
) lut_6_10 (
    .O(x6_y10),
    .I0(x4_y12),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110111000110)
) lut_7_10 (
    .O(x7_y10),
    .I0(x4_y13),
    .I1(x5_y13),
    .I2(x5_y8),
    .I3(x5_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111001100011)
) lut_8_10 (
    .O(x8_y10),
    .I0(x6_y14),
    .I1(1'b0),
    .I2(x5_y11),
    .I3(x5_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111000110000)
) lut_9_10 (
    .O(x9_y10),
    .I0(x7_y14),
    .I1(1'b0),
    .I2(x5_y11),
    .I3(x5_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111011010111)
) lut_10_10 (
    .O(x10_y10),
    .I0(x8_y11),
    .I1(x8_y7),
    .I2(1'b0),
    .I3(x7_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010101101101)
) lut_11_10 (
    .O(x11_y10),
    .I0(x9_y10),
    .I1(x9_y12),
    .I2(x9_y7),
    .I3(x9_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010011001101)
) lut_12_10 (
    .O(x12_y10),
    .I0(1'b0),
    .I1(x10_y8),
    .I2(x9_y7),
    .I3(x9_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101011000011)
) lut_13_10 (
    .O(x13_y10),
    .I0(x10_y8),
    .I1(x11_y14),
    .I2(x10_y5),
    .I3(x11_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100001101101)
) lut_14_10 (
    .O(x14_y10),
    .I0(x12_y11),
    .I1(1'b0),
    .I2(x11_y6),
    .I3(x12_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100011011011)
) lut_15_10 (
    .O(x15_y10),
    .I0(x13_y9),
    .I1(x13_y13),
    .I2(x12_y10),
    .I3(x13_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010110010010)
) lut_16_10 (
    .O(x16_y10),
    .I0(1'b0),
    .I1(x14_y15),
    .I2(x13_y8),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110011000001)
) lut_17_10 (
    .O(x17_y10),
    .I0(1'b0),
    .I1(x15_y9),
    .I2(x14_y13),
    .I3(x14_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111101111001)
) lut_18_10 (
    .O(x18_y10),
    .I0(x16_y8),
    .I1(x16_y5),
    .I2(x15_y10),
    .I3(x16_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010000010101)
) lut_19_10 (
    .O(x19_y10),
    .I0(x17_y9),
    .I1(x16_y9),
    .I2(x16_y8),
    .I3(x16_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100001110011)
) lut_20_10 (
    .O(x20_y10),
    .I0(1'b0),
    .I1(x18_y6),
    .I2(x18_y7),
    .I3(x17_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111111000001)
) lut_21_10 (
    .O(x21_y10),
    .I0(x19_y5),
    .I1(1'b0),
    .I2(x18_y5),
    .I3(x19_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100001110011)
) lut_22_10 (
    .O(x22_y10),
    .I0(x19_y13),
    .I1(x20_y10),
    .I2(x19_y10),
    .I3(x20_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001001100001)
) lut_23_10 (
    .O(x23_y10),
    .I0(x20_y6),
    .I1(x21_y6),
    .I2(x20_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010110011000)
) lut_24_10 (
    .O(x24_y10),
    .I0(x22_y15),
    .I1(x21_y14),
    .I2(x22_y13),
    .I3(x21_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111010111110)
) lut_25_10 (
    .O(x25_y10),
    .I0(x23_y11),
    .I1(x23_y12),
    .I2(x23_y10),
    .I3(x22_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001101010001)
) lut_26_10 (
    .O(x26_y10),
    .I0(x24_y5),
    .I1(x24_y6),
    .I2(x24_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000000001011)
) lut_27_10 (
    .O(x27_y10),
    .I0(x25_y6),
    .I1(x24_y5),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011010100011)
) lut_28_10 (
    .O(x28_y10),
    .I0(1'b0),
    .I1(x26_y7),
    .I2(x25_y13),
    .I3(x25_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000001011110)
) lut_29_10 (
    .O(x29_y10),
    .I0(1'b0),
    .I1(x27_y8),
    .I2(x26_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100000101111)
) lut_30_10 (
    .O(x30_y10),
    .I0(x28_y13),
    .I1(x28_y5),
    .I2(x28_y15),
    .I3(x27_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100010101101)
) lut_31_10 (
    .O(x31_y10),
    .I0(x29_y11),
    .I1(1'b0),
    .I2(x29_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000001110011)
) lut_32_10 (
    .O(x32_y10),
    .I0(x30_y9),
    .I1(x29_y11),
    .I2(x30_y8),
    .I3(x29_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100101101111)
) lut_33_10 (
    .O(x33_y10),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x31_y11),
    .I3(x31_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010010101000)
) lut_34_10 (
    .O(x34_y10),
    .I0(x32_y5),
    .I1(x31_y9),
    .I2(x31_y12),
    .I3(x31_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110100101110)
) lut_35_10 (
    .O(x35_y10),
    .I0(1'b0),
    .I1(x32_y6),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011010000100)
) lut_36_10 (
    .O(x36_y10),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x33_y14),
    .I3(x34_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101100010111)
) lut_37_10 (
    .O(x37_y10),
    .I0(1'b0),
    .I1(x34_y9),
    .I2(x35_y9),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011100111011)
) lut_38_10 (
    .O(x38_y10),
    .I0(x36_y10),
    .I1(x36_y12),
    .I2(x36_y9),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010101010100)
) lut_39_10 (
    .O(x39_y10),
    .I0(x36_y10),
    .I1(x36_y6),
    .I2(x37_y8),
    .I3(x36_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101110101101)
) lut_40_10 (
    .O(x40_y10),
    .I0(1'b0),
    .I1(x37_y14),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011001111010)
) lut_41_10 (
    .O(x41_y10),
    .I0(x38_y8),
    .I1(x39_y6),
    .I2(x38_y7),
    .I3(x39_y5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100101001110)
) lut_42_10 (
    .O(x42_y10),
    .I0(x40_y14),
    .I1(x40_y5),
    .I2(x39_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101000010001)
) lut_43_10 (
    .O(x43_y10),
    .I0(x41_y8),
    .I1(x40_y11),
    .I2(x40_y13),
    .I3(x40_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011110100100)
) lut_44_10 (
    .O(x44_y10),
    .I0(x41_y5),
    .I1(x41_y8),
    .I2(x42_y14),
    .I3(x41_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110101101101)
) lut_45_10 (
    .O(x45_y10),
    .I0(x43_y10),
    .I1(x42_y10),
    .I2(x42_y8),
    .I3(x42_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100010011101)
) lut_46_10 (
    .O(x46_y10),
    .I0(x44_y11),
    .I1(1'b0),
    .I2(x44_y10),
    .I3(x43_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001011000010)
) lut_47_10 (
    .O(x47_y10),
    .I0(x45_y15),
    .I1(x45_y14),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101111001111)
) lut_48_10 (
    .O(x48_y10),
    .I0(x45_y9),
    .I1(x46_y13),
    .I2(x46_y11),
    .I3(x45_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010101101110)
) lut_49_10 (
    .O(x49_y10),
    .I0(x46_y12),
    .I1(1'b0),
    .I2(x47_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000000001110)
) lut_50_10 (
    .O(x50_y10),
    .I0(1'b0),
    .I1(x48_y14),
    .I2(x47_y7),
    .I3(x47_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001011110110)
) lut_51_10 (
    .O(x51_y10),
    .I0(x49_y14),
    .I1(x49_y5),
    .I2(x49_y9),
    .I3(x48_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011000000011)
) lut_52_10 (
    .O(x52_y10),
    .I0(x49_y13),
    .I1(x49_y5),
    .I2(x50_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001001001010)
) lut_53_10 (
    .O(x53_y10),
    .I0(x50_y8),
    .I1(x50_y13),
    .I2(1'b0),
    .I3(x51_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011110100110)
) lut_54_10 (
    .O(x54_y10),
    .I0(x51_y7),
    .I1(x52_y6),
    .I2(x51_y9),
    .I3(x52_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010010001100)
) lut_55_10 (
    .O(x55_y10),
    .I0(x52_y11),
    .I1(x53_y12),
    .I2(x52_y15),
    .I3(x52_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110010110001)
) lut_56_10 (
    .O(x56_y10),
    .I0(x54_y9),
    .I1(x54_y6),
    .I2(1'b0),
    .I3(x53_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100011000000)
) lut_57_10 (
    .O(x57_y10),
    .I0(x54_y14),
    .I1(x54_y13),
    .I2(x54_y5),
    .I3(x54_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000010000100)
) lut_58_10 (
    .O(x58_y10),
    .I0(x55_y5),
    .I1(x56_y14),
    .I2(x55_y10),
    .I3(x55_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011001101110)
) lut_59_10 (
    .O(x59_y10),
    .I0(x57_y5),
    .I1(x56_y11),
    .I2(x56_y12),
    .I3(x57_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101110010100)
) lut_60_10 (
    .O(x60_y10),
    .I0(1'b0),
    .I1(x57_y8),
    .I2(1'b0),
    .I3(x58_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111010001101)
) lut_61_10 (
    .O(x61_y10),
    .I0(x58_y13),
    .I1(1'b0),
    .I2(x59_y12),
    .I3(x59_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011010010110)
) lut_62_10 (
    .O(x62_y10),
    .I0(x59_y12),
    .I1(x60_y7),
    .I2(x59_y8),
    .I3(x60_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110000000010)
) lut_0_11 (
    .O(x0_y11),
    .I0(1'b0),
    .I1(in1),
    .I2(in7),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010001101001)
) lut_1_11 (
    .O(x1_y11),
    .I0(in0),
    .I1(in6),
    .I2(in9),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000110111001)
) lut_2_11 (
    .O(x2_y11),
    .I0(1'b0),
    .I1(1'b0),
    .I2(in1),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110001100011)
) lut_3_11 (
    .O(x3_y11),
    .I0(1'b0),
    .I1(in6),
    .I2(x1_y15),
    .I3(x1_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101010000000)
) lut_4_11 (
    .O(x4_y11),
    .I0(1'b0),
    .I1(x2_y16),
    .I2(1'b0),
    .I3(x1_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011010000111)
) lut_5_11 (
    .O(x5_y11),
    .I0(x3_y14),
    .I1(x2_y12),
    .I2(x3_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001110100000)
) lut_6_11 (
    .O(x6_y11),
    .I0(x3_y15),
    .I1(1'b0),
    .I2(x4_y15),
    .I3(x3_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110001101001)
) lut_7_11 (
    .O(x7_y11),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x4_y16),
    .I3(x4_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100011011010)
) lut_8_11 (
    .O(x8_y11),
    .I0(x5_y11),
    .I1(x6_y10),
    .I2(x5_y14),
    .I3(x5_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110110110010)
) lut_9_11 (
    .O(x9_y11),
    .I0(x7_y6),
    .I1(x7_y15),
    .I2(x5_y14),
    .I3(x5_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000011010011)
) lut_10_11 (
    .O(x10_y11),
    .I0(x7_y16),
    .I1(x7_y9),
    .I2(x8_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101001010111)
) lut_11_11 (
    .O(x11_y11),
    .I0(x9_y7),
    .I1(x8_y16),
    .I2(x9_y8),
    .I3(x9_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011001110101)
) lut_12_11 (
    .O(x12_y11),
    .I0(x10_y8),
    .I1(x9_y10),
    .I2(x9_y15),
    .I3(x9_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110000000111)
) lut_13_11 (
    .O(x13_y11),
    .I0(x11_y11),
    .I1(x10_y11),
    .I2(x10_y16),
    .I3(x10_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111110001111)
) lut_14_11 (
    .O(x14_y11),
    .I0(x12_y13),
    .I1(x12_y15),
    .I2(1'b0),
    .I3(x11_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111010110010)
) lut_15_11 (
    .O(x15_y11),
    .I0(x13_y13),
    .I1(1'b0),
    .I2(x13_y8),
    .I3(x13_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001100101011)
) lut_16_11 (
    .O(x16_y11),
    .I0(x13_y16),
    .I1(x13_y14),
    .I2(x13_y8),
    .I3(x13_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110001001101)
) lut_17_11 (
    .O(x17_y11),
    .I0(x14_y16),
    .I1(x14_y6),
    .I2(x14_y7),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001000101110)
) lut_18_11 (
    .O(x18_y11),
    .I0(x15_y13),
    .I1(x15_y12),
    .I2(x15_y12),
    .I3(x16_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011110001000)
) lut_19_11 (
    .O(x19_y11),
    .I0(x17_y6),
    .I1(x17_y8),
    .I2(x16_y11),
    .I3(x17_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001001110001)
) lut_20_11 (
    .O(x20_y11),
    .I0(x18_y10),
    .I1(x17_y14),
    .I2(x17_y8),
    .I3(x17_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000010111101)
) lut_21_11 (
    .O(x21_y11),
    .I0(x19_y14),
    .I1(x18_y7),
    .I2(x19_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100111110011)
) lut_22_11 (
    .O(x22_y11),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x19_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000010110000)
) lut_23_11 (
    .O(x23_y11),
    .I0(x21_y8),
    .I1(x20_y12),
    .I2(x21_y12),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010101001111)
) lut_24_11 (
    .O(x24_y11),
    .I0(x21_y13),
    .I1(x21_y15),
    .I2(x22_y15),
    .I3(x21_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000001101110)
) lut_25_11 (
    .O(x25_y11),
    .I0(x23_y16),
    .I1(x22_y15),
    .I2(x23_y12),
    .I3(x22_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000011110011)
) lut_26_11 (
    .O(x26_y11),
    .I0(x24_y16),
    .I1(x23_y9),
    .I2(x23_y16),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011001100101)
) lut_27_11 (
    .O(x27_y11),
    .I0(1'b0),
    .I1(x24_y10),
    .I2(1'b0),
    .I3(x24_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101001000001)
) lut_28_11 (
    .O(x28_y11),
    .I0(x26_y8),
    .I1(x26_y12),
    .I2(x26_y10),
    .I3(x25_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000110111001)
) lut_29_11 (
    .O(x29_y11),
    .I0(x26_y14),
    .I1(x27_y13),
    .I2(1'b0),
    .I3(x27_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100101001101)
) lut_30_11 (
    .O(x30_y11),
    .I0(x27_y14),
    .I1(x28_y8),
    .I2(1'b0),
    .I3(x28_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110100001100)
) lut_31_11 (
    .O(x31_y11),
    .I0(1'b0),
    .I1(x29_y7),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011100111010)
) lut_32_11 (
    .O(x32_y11),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x30_y7),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000001010001)
) lut_33_11 (
    .O(x33_y11),
    .I0(x30_y10),
    .I1(x31_y10),
    .I2(x30_y12),
    .I3(x30_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110000010011)
) lut_34_11 (
    .O(x34_y11),
    .I0(x31_y13),
    .I1(x32_y14),
    .I2(1'b0),
    .I3(x31_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000010100001)
) lut_35_11 (
    .O(x35_y11),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x32_y7),
    .I3(x32_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000110111010)
) lut_36_11 (
    .O(x36_y11),
    .I0(x33_y12),
    .I1(x33_y9),
    .I2(x34_y11),
    .I3(x34_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101000101011)
) lut_37_11 (
    .O(x37_y11),
    .I0(1'b0),
    .I1(x34_y14),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100010110110)
) lut_38_11 (
    .O(x38_y11),
    .I0(1'b0),
    .I1(x36_y12),
    .I2(x35_y15),
    .I3(x36_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001010010010)
) lut_39_11 (
    .O(x39_y11),
    .I0(x36_y11),
    .I1(x37_y11),
    .I2(x36_y10),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001101110110)
) lut_40_11 (
    .O(x40_y11),
    .I0(x38_y6),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x37_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111101000000)
) lut_41_11 (
    .O(x41_y11),
    .I0(x38_y14),
    .I1(x38_y15),
    .I2(x39_y12),
    .I3(x38_y6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000111000011)
) lut_42_11 (
    .O(x42_y11),
    .I0(x40_y11),
    .I1(x40_y16),
    .I2(x40_y7),
    .I3(x40_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010100011110)
) lut_43_11 (
    .O(x43_y11),
    .I0(x40_y15),
    .I1(x40_y15),
    .I2(x40_y12),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111010010111)
) lut_44_11 (
    .O(x44_y11),
    .I0(x42_y11),
    .I1(x41_y12),
    .I2(1'b0),
    .I3(x41_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111010101101)
) lut_45_11 (
    .O(x45_y11),
    .I0(x43_y10),
    .I1(1'b0),
    .I2(x42_y9),
    .I3(x43_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001111111000)
) lut_46_11 (
    .O(x46_y11),
    .I0(x43_y10),
    .I1(x44_y14),
    .I2(x43_y9),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000101000100)
) lut_47_11 (
    .O(x47_y11),
    .I0(x44_y15),
    .I1(x45_y10),
    .I2(x45_y12),
    .I3(x45_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001110101100)
) lut_48_11 (
    .O(x48_y11),
    .I0(x46_y9),
    .I1(x45_y9),
    .I2(x45_y11),
    .I3(x45_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100100100010)
) lut_49_11 (
    .O(x49_y11),
    .I0(1'b0),
    .I1(x46_y7),
    .I2(x46_y10),
    .I3(x46_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010001110011)
) lut_50_11 (
    .O(x50_y11),
    .I0(1'b0),
    .I1(x48_y11),
    .I2(x47_y12),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001111011110)
) lut_51_11 (
    .O(x51_y11),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x48_y9),
    .I3(x48_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101100010011)
) lut_52_11 (
    .O(x52_y11),
    .I0(x50_y8),
    .I1(1'b0),
    .I2(x50_y7),
    .I3(x49_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111011011110)
) lut_53_11 (
    .O(x53_y11),
    .I0(x51_y8),
    .I1(x50_y15),
    .I2(x51_y14),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111011101100)
) lut_54_11 (
    .O(x54_y11),
    .I0(x51_y10),
    .I1(1'b0),
    .I2(x51_y6),
    .I3(x51_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010101111110)
) lut_55_11 (
    .O(x55_y11),
    .I0(1'b0),
    .I1(x53_y15),
    .I2(x53_y15),
    .I3(x53_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100000101001)
) lut_56_11 (
    .O(x56_y11),
    .I0(x53_y6),
    .I1(x54_y11),
    .I2(x53_y14),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000000010111)
) lut_57_11 (
    .O(x57_y11),
    .I0(x54_y6),
    .I1(x54_y15),
    .I2(x55_y16),
    .I3(x55_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100100101100)
) lut_58_11 (
    .O(x58_y11),
    .I0(1'b0),
    .I1(x56_y16),
    .I2(1'b0),
    .I3(x56_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010010011011)
) lut_59_11 (
    .O(x59_y11),
    .I0(x56_y16),
    .I1(x57_y12),
    .I2(1'b0),
    .I3(x56_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001001000011)
) lut_60_11 (
    .O(x60_y11),
    .I0(x57_y13),
    .I1(1'b0),
    .I2(x57_y10),
    .I3(x58_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010110110000)
) lut_61_11 (
    .O(x61_y11),
    .I0(x58_y14),
    .I1(x59_y12),
    .I2(1'b0),
    .I3(x58_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001101110101)
) lut_62_11 (
    .O(x62_y11),
    .I0(x60_y7),
    .I1(x59_y8),
    .I2(x59_y9),
    .I3(x60_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011110010100)
) lut_0_12 (
    .O(x0_y12),
    .I0(in7),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111000101111)
) lut_1_12 (
    .O(x1_y12),
    .I0(1'b0),
    .I1(in5),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110000000000)
) lut_2_12 (
    .O(x2_y12),
    .I0(in7),
    .I1(in4),
    .I2(1'b0),
    .I3(in7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000001110010)
) lut_3_12 (
    .O(x3_y12),
    .I0(in9),
    .I1(x1_y17),
    .I2(in4),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010001111111)
) lut_4_12 (
    .O(x4_y12),
    .I0(x1_y15),
    .I1(x1_y7),
    .I2(1'b0),
    .I3(x1_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001011100001)
) lut_5_12 (
    .O(x5_y12),
    .I0(1'b0),
    .I1(x2_y8),
    .I2(1'b0),
    .I3(x2_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100010010010)
) lut_6_12 (
    .O(x6_y12),
    .I0(1'b0),
    .I1(x4_y11),
    .I2(x3_y9),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101100011010)
) lut_7_12 (
    .O(x7_y12),
    .I0(x4_y12),
    .I1(x4_y13),
    .I2(x5_y12),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011100010100)
) lut_8_12 (
    .O(x8_y12),
    .I0(x5_y17),
    .I1(x5_y8),
    .I2(x6_y9),
    .I3(x6_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110011000010)
) lut_9_12 (
    .O(x9_y12),
    .I0(x6_y12),
    .I1(x6_y11),
    .I2(x6_y9),
    .I3(x6_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111010110001)
) lut_10_12 (
    .O(x10_y12),
    .I0(x8_y7),
    .I1(1'b0),
    .I2(x7_y10),
    .I3(x7_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010100110100)
) lut_11_12 (
    .O(x11_y12),
    .I0(x9_y15),
    .I1(x8_y17),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111100000101)
) lut_12_12 (
    .O(x12_y12),
    .I0(x9_y14),
    .I1(x10_y11),
    .I2(x9_y13),
    .I3(x10_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111110000110)
) lut_13_12 (
    .O(x13_y12),
    .I0(x10_y9),
    .I1(x10_y10),
    .I2(x11_y17),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100011111011)
) lut_14_12 (
    .O(x14_y12),
    .I0(x12_y13),
    .I1(x11_y12),
    .I2(x12_y12),
    .I3(x12_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110100001011)
) lut_15_12 (
    .O(x15_y12),
    .I0(x13_y11),
    .I1(x13_y7),
    .I2(x12_y16),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110011101001)
) lut_16_12 (
    .O(x16_y12),
    .I0(1'b0),
    .I1(x14_y11),
    .I2(x13_y15),
    .I3(x13_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000010110010)
) lut_17_12 (
    .O(x17_y12),
    .I0(x15_y14),
    .I1(x15_y13),
    .I2(x14_y16),
    .I3(x15_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000001101011)
) lut_18_12 (
    .O(x18_y12),
    .I0(x15_y14),
    .I1(x15_y10),
    .I2(1'b0),
    .I3(x16_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010000000101)
) lut_19_12 (
    .O(x19_y12),
    .I0(x16_y14),
    .I1(x16_y13),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001001011011)
) lut_20_12 (
    .O(x20_y12),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x17_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110011110010)
) lut_21_12 (
    .O(x21_y12),
    .I0(x18_y17),
    .I1(1'b0),
    .I2(x18_y16),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101000010011)
) lut_22_12 (
    .O(x22_y12),
    .I0(x19_y9),
    .I1(1'b0),
    .I2(x19_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111100101111)
) lut_23_12 (
    .O(x23_y12),
    .I0(x21_y8),
    .I1(x21_y12),
    .I2(1'b0),
    .I3(x21_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011100010010)
) lut_24_12 (
    .O(x24_y12),
    .I0(x22_y8),
    .I1(x22_y7),
    .I2(x21_y9),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001011111100)
) lut_25_12 (
    .O(x25_y12),
    .I0(x22_y16),
    .I1(x22_y15),
    .I2(1'b0),
    .I3(x22_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110001111011)
) lut_26_12 (
    .O(x26_y12),
    .I0(x23_y11),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x23_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111110110011)
) lut_27_12 (
    .O(x27_y12),
    .I0(x24_y12),
    .I1(x24_y13),
    .I2(1'b0),
    .I3(x25_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011101111011)
) lut_28_12 (
    .O(x28_y12),
    .I0(x26_y12),
    .I1(x26_y12),
    .I2(x25_y16),
    .I3(x25_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011001000110)
) lut_29_12 (
    .O(x29_y12),
    .I0(x26_y10),
    .I1(x27_y15),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111000100100)
) lut_30_12 (
    .O(x30_y12),
    .I0(x27_y9),
    .I1(x27_y11),
    .I2(1'b0),
    .I3(x28_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010101010110)
) lut_31_12 (
    .O(x31_y12),
    .I0(x28_y10),
    .I1(x28_y13),
    .I2(x29_y14),
    .I3(x28_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101101110001)
) lut_32_12 (
    .O(x32_y12),
    .I0(x30_y11),
    .I1(x29_y11),
    .I2(x29_y7),
    .I3(x30_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110110110011)
) lut_33_12 (
    .O(x33_y12),
    .I0(x30_y16),
    .I1(1'b0),
    .I2(x30_y13),
    .I3(x31_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111010010101)
) lut_34_12 (
    .O(x34_y12),
    .I0(x32_y7),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x31_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101001010000)
) lut_35_12 (
    .O(x35_y12),
    .I0(x33_y15),
    .I1(1'b0),
    .I2(x32_y7),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111011100110)
) lut_36_12 (
    .O(x36_y12),
    .I0(x34_y17),
    .I1(x34_y17),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110110101100)
) lut_37_12 (
    .O(x37_y12),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x34_y14),
    .I3(x34_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111100100000)
) lut_38_12 (
    .O(x38_y12),
    .I0(x36_y13),
    .I1(x35_y12),
    .I2(1'b0),
    .I3(x36_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101100000100)
) lut_39_12 (
    .O(x39_y12),
    .I0(x36_y16),
    .I1(x36_y16),
    .I2(1'b0),
    .I3(x37_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100000110011)
) lut_40_12 (
    .O(x40_y12),
    .I0(x38_y17),
    .I1(x38_y13),
    .I2(x38_y15),
    .I3(x38_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000000000011)
) lut_41_12 (
    .O(x41_y12),
    .I0(x39_y13),
    .I1(x39_y10),
    .I2(1'b0),
    .I3(x39_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101111011000)
) lut_42_12 (
    .O(x42_y12),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x40_y13),
    .I3(x39_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100111101001)
) lut_43_12 (
    .O(x43_y12),
    .I0(x41_y7),
    .I1(x41_y14),
    .I2(1'b0),
    .I3(x41_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110010101001)
) lut_44_12 (
    .O(x44_y12),
    .I0(x41_y15),
    .I1(1'b0),
    .I2(x42_y12),
    .I3(x42_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001101011111)
) lut_45_12 (
    .O(x45_y12),
    .I0(x43_y15),
    .I1(x43_y17),
    .I2(x42_y16),
    .I3(x42_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111110010110)
) lut_46_12 (
    .O(x46_y12),
    .I0(x43_y17),
    .I1(x43_y13),
    .I2(x43_y11),
    .I3(x43_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101100011111)
) lut_47_12 (
    .O(x47_y12),
    .I0(x45_y12),
    .I1(x44_y10),
    .I2(1'b0),
    .I3(x44_y7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111000110101)
) lut_48_12 (
    .O(x48_y12),
    .I0(x46_y7),
    .I1(x45_y12),
    .I2(x45_y14),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100101010101)
) lut_49_12 (
    .O(x49_y12),
    .I0(x46_y12),
    .I1(x47_y9),
    .I2(x46_y7),
    .I3(x46_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001100100110)
) lut_50_12 (
    .O(x50_y12),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x48_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101111100110)
) lut_51_12 (
    .O(x51_y12),
    .I0(1'b0),
    .I1(x48_y7),
    .I2(x49_y10),
    .I3(x49_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110000110010)
) lut_52_12 (
    .O(x52_y12),
    .I0(x50_y17),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x49_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001010101000)
) lut_53_12 (
    .O(x53_y12),
    .I0(x51_y12),
    .I1(x50_y11),
    .I2(x51_y10),
    .I3(x50_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011111010010)
) lut_54_12 (
    .O(x54_y12),
    .I0(x51_y12),
    .I1(x52_y13),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011110100111)
) lut_55_12 (
    .O(x55_y12),
    .I0(1'b0),
    .I1(x53_y14),
    .I2(x52_y14),
    .I3(x53_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111011101110)
) lut_56_12 (
    .O(x56_y12),
    .I0(x54_y11),
    .I1(x54_y7),
    .I2(x54_y9),
    .I3(x53_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011101010000)
) lut_57_12 (
    .O(x57_y12),
    .I0(x55_y16),
    .I1(x54_y14),
    .I2(x55_y10),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010011111000)
) lut_58_12 (
    .O(x58_y12),
    .I0(x56_y11),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x56_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010001010010)
) lut_59_12 (
    .O(x59_y12),
    .I0(1'b0),
    .I1(x57_y14),
    .I2(x56_y14),
    .I3(x56_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110011110101)
) lut_60_12 (
    .O(x60_y12),
    .I0(1'b0),
    .I1(x57_y9),
    .I2(x57_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111001101100)
) lut_61_12 (
    .O(x61_y12),
    .I0(x58_y12),
    .I1(x58_y16),
    .I2(x58_y10),
    .I3(x59_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001110110110)
) lut_62_12 (
    .O(x62_y12),
    .I0(1'b0),
    .I1(x59_y15),
    .I2(x59_y17),
    .I3(x60_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010001011010)
) lut_0_13 (
    .O(x0_y13),
    .I0(in7),
    .I1(1'b0),
    .I2(1'b0),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111110100100)
) lut_1_13 (
    .O(x1_y13),
    .I0(in9),
    .I1(in3),
    .I2(in3),
    .I3(in3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010010100101)
) lut_2_13 (
    .O(x2_y13),
    .I0(in7),
    .I1(1'b0),
    .I2(in3),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001000010100)
) lut_3_13 (
    .O(x3_y13),
    .I0(in0),
    .I1(1'b0),
    .I2(in7),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101011010111)
) lut_4_13 (
    .O(x4_y13),
    .I0(x1_y15),
    .I1(x1_y17),
    .I2(x2_y15),
    .I3(x1_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111011110011)
) lut_5_13 (
    .O(x5_y13),
    .I0(1'b0),
    .I1(x3_y16),
    .I2(x2_y15),
    .I3(x3_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100000001000)
) lut_6_13 (
    .O(x6_y13),
    .I0(x3_y15),
    .I1(x3_y8),
    .I2(x3_y17),
    .I3(x4_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010110101100)
) lut_7_13 (
    .O(x7_y13),
    .I0(x4_y9),
    .I1(x5_y18),
    .I2(x4_y10),
    .I3(x5_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000100001111)
) lut_8_13 (
    .O(x8_y13),
    .I0(1'b0),
    .I1(x6_y17),
    .I2(x5_y18),
    .I3(x5_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010111000010)
) lut_9_13 (
    .O(x9_y13),
    .I0(x6_y17),
    .I1(x7_y18),
    .I2(x5_y18),
    .I3(x5_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011100110000)
) lut_10_13 (
    .O(x10_y13),
    .I0(x8_y18),
    .I1(x8_y11),
    .I2(1'b0),
    .I3(x8_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101011110001)
) lut_11_13 (
    .O(x11_y13),
    .I0(1'b0),
    .I1(x8_y15),
    .I2(1'b0),
    .I3(x8_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010110011000)
) lut_12_13 (
    .O(x12_y13),
    .I0(1'b0),
    .I1(x10_y15),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001011001010)
) lut_13_13 (
    .O(x13_y13),
    .I0(x10_y16),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x11_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001010001110)
) lut_14_13 (
    .O(x14_y13),
    .I0(x12_y11),
    .I1(x11_y11),
    .I2(x12_y9),
    .I3(x11_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000000100100)
) lut_15_13 (
    .O(x15_y13),
    .I0(x13_y17),
    .I1(x12_y15),
    .I2(x13_y13),
    .I3(x13_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110011001001)
) lut_16_13 (
    .O(x16_y13),
    .I0(1'b0),
    .I1(x14_y15),
    .I2(x14_y10),
    .I3(x14_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110010101111)
) lut_17_13 (
    .O(x17_y13),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x15_y16),
    .I3(x14_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010100011101)
) lut_18_13 (
    .O(x18_y13),
    .I0(x16_y10),
    .I1(x15_y10),
    .I2(x16_y16),
    .I3(x15_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001100101110)
) lut_19_13 (
    .O(x19_y13),
    .I0(x17_y18),
    .I1(x17_y16),
    .I2(1'b0),
    .I3(x16_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101111011101)
) lut_20_13 (
    .O(x20_y13),
    .I0(1'b0),
    .I1(x17_y11),
    .I2(x17_y17),
    .I3(x17_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010100110011)
) lut_21_13 (
    .O(x21_y13),
    .I0(x18_y15),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101101000111)
) lut_22_13 (
    .O(x22_y13),
    .I0(x20_y9),
    .I1(1'b0),
    .I2(x20_y8),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000100110001)
) lut_23_13 (
    .O(x23_y13),
    .I0(x20_y12),
    .I1(x20_y10),
    .I2(1'b0),
    .I3(x21_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110011101001)
) lut_24_13 (
    .O(x24_y13),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x21_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001101001010)
) lut_25_13 (
    .O(x25_y13),
    .I0(x23_y17),
    .I1(1'b0),
    .I2(x22_y15),
    .I3(x23_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001110101001)
) lut_26_13 (
    .O(x26_y13),
    .I0(1'b0),
    .I1(x23_y16),
    .I2(1'b0),
    .I3(x24_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100011001001)
) lut_27_13 (
    .O(x27_y13),
    .I0(x25_y16),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x25_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001000111110)
) lut_28_13 (
    .O(x28_y13),
    .I0(x26_y14),
    .I1(x25_y18),
    .I2(1'b0),
    .I3(x26_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101010011001)
) lut_29_13 (
    .O(x29_y13),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x26_y9),
    .I3(x26_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101110010001)
) lut_30_13 (
    .O(x30_y13),
    .I0(x27_y11),
    .I1(x27_y13),
    .I2(x27_y11),
    .I3(x28_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101000000110)
) lut_31_13 (
    .O(x31_y13),
    .I0(x29_y15),
    .I1(x29_y10),
    .I2(1'b0),
    .I3(x28_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010001010001)
) lut_32_13 (
    .O(x32_y13),
    .I0(x30_y9),
    .I1(x29_y18),
    .I2(x30_y9),
    .I3(x30_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001101101111)
) lut_33_13 (
    .O(x33_y13),
    .I0(1'b0),
    .I1(x31_y15),
    .I2(x31_y17),
    .I3(x31_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110111011011)
) lut_34_13 (
    .O(x34_y13),
    .I0(x31_y8),
    .I1(x32_y11),
    .I2(x32_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100000000010)
) lut_35_13 (
    .O(x35_y13),
    .I0(1'b0),
    .I1(x32_y12),
    .I2(x33_y9),
    .I3(x32_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100110101010)
) lut_36_13 (
    .O(x36_y13),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x33_y12),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011001010001)
) lut_37_13 (
    .O(x37_y13),
    .I0(x34_y10),
    .I1(x35_y13),
    .I2(x35_y14),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111111111001)
) lut_38_13 (
    .O(x38_y13),
    .I0(x35_y17),
    .I1(1'b0),
    .I2(x35_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011010111010)
) lut_39_13 (
    .O(x39_y13),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x36_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111010011111)
) lut_40_13 (
    .O(x40_y13),
    .I0(x37_y14),
    .I1(x38_y14),
    .I2(x37_y11),
    .I3(x38_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101000110100)
) lut_41_13 (
    .O(x41_y13),
    .I0(x39_y15),
    .I1(1'b0),
    .I2(x39_y11),
    .I3(x39_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110010000101)
) lut_42_13 (
    .O(x42_y13),
    .I0(x39_y16),
    .I1(x40_y13),
    .I2(x39_y13),
    .I3(x40_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000011100000)
) lut_43_13 (
    .O(x43_y13),
    .I0(x40_y9),
    .I1(x40_y17),
    .I2(x41_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110110011101)
) lut_44_13 (
    .O(x44_y13),
    .I0(1'b0),
    .I1(x42_y15),
    .I2(x41_y9),
    .I3(x42_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101000010000)
) lut_45_13 (
    .O(x45_y13),
    .I0(1'b0),
    .I1(x42_y16),
    .I2(1'b0),
    .I3(x43_y8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010001101100)
) lut_46_13 (
    .O(x46_y13),
    .I0(x44_y13),
    .I1(1'b0),
    .I2(x44_y16),
    .I3(x43_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010101100011)
) lut_47_13 (
    .O(x47_y13),
    .I0(x44_y18),
    .I1(x45_y15),
    .I2(1'b0),
    .I3(x44_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011101000000)
) lut_48_13 (
    .O(x48_y13),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x46_y10),
    .I3(x46_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111111001000)
) lut_49_13 (
    .O(x49_y13),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x46_y10),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010111001111)
) lut_50_13 (
    .O(x50_y13),
    .I0(x48_y8),
    .I1(1'b0),
    .I2(x48_y13),
    .I3(x47_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000010110000)
) lut_51_13 (
    .O(x51_y13),
    .I0(x48_y9),
    .I1(x48_y9),
    .I2(x49_y16),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101101110001)
) lut_52_13 (
    .O(x52_y13),
    .I0(x50_y8),
    .I1(x50_y9),
    .I2(x50_y12),
    .I3(x50_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110000101100)
) lut_53_13 (
    .O(x53_y13),
    .I0(x51_y18),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x51_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100010111110)
) lut_54_13 (
    .O(x54_y13),
    .I0(x52_y8),
    .I1(1'b0),
    .I2(x52_y17),
    .I3(x52_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011011010010)
) lut_55_13 (
    .O(x55_y13),
    .I0(x53_y8),
    .I1(x52_y13),
    .I2(x53_y15),
    .I3(x53_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000100011111)
) lut_56_13 (
    .O(x56_y13),
    .I0(x54_y9),
    .I1(x53_y14),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110100111011)
) lut_57_13 (
    .O(x57_y13),
    .I0(x55_y9),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x55_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000110000110)
) lut_58_13 (
    .O(x58_y13),
    .I0(x55_y17),
    .I1(x55_y13),
    .I2(x56_y8),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001010101101)
) lut_59_13 (
    .O(x59_y13),
    .I0(x56_y9),
    .I1(x56_y18),
    .I2(x57_y12),
    .I3(x57_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011011010111)
) lut_60_13 (
    .O(x60_y13),
    .I0(x57_y12),
    .I1(x58_y16),
    .I2(x58_y13),
    .I3(x58_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111101000010)
) lut_61_13 (
    .O(x61_y13),
    .I0(x58_y17),
    .I1(x59_y8),
    .I2(x59_y17),
    .I3(x59_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001010101101)
) lut_62_13 (
    .O(x62_y13),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x60_y10),
    .I3(x60_y9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100000000001)
) lut_0_14 (
    .O(x0_y14),
    .I0(in6),
    .I1(in6),
    .I2(in4),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100010101110)
) lut_1_14 (
    .O(x1_y14),
    .I0(in1),
    .I1(in2),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111010010101)
) lut_2_14 (
    .O(x2_y14),
    .I0(in3),
    .I1(in8),
    .I2(in0),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110111100111)
) lut_3_14 (
    .O(x3_y14),
    .I0(x1_y17),
    .I1(in1),
    .I2(1'b0),
    .I3(x1_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100000000000)
) lut_4_14 (
    .O(x4_y14),
    .I0(x2_y16),
    .I1(1'b0),
    .I2(x1_y16),
    .I3(x2_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001011010111)
) lut_5_14 (
    .O(x5_y14),
    .I0(x3_y9),
    .I1(x2_y15),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111011011001)
) lut_6_14 (
    .O(x6_y14),
    .I0(x3_y10),
    .I1(1'b0),
    .I2(x3_y15),
    .I3(x4_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110101111110)
) lut_7_14 (
    .O(x7_y14),
    .I0(x4_y10),
    .I1(x4_y12),
    .I2(1'b0),
    .I3(x4_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100001010010)
) lut_8_14 (
    .O(x8_y14),
    .I0(x5_y11),
    .I1(x5_y16),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100001100101)
) lut_9_14 (
    .O(x9_y14),
    .I0(x7_y13),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100100100011)
) lut_10_14 (
    .O(x10_y14),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x7_y16),
    .I3(x8_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100011001001)
) lut_11_14 (
    .O(x11_y14),
    .I0(x8_y19),
    .I1(x8_y9),
    .I2(x8_y16),
    .I3(x8_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101000001000)
) lut_12_14 (
    .O(x12_y14),
    .I0(x9_y13),
    .I1(x10_y18),
    .I2(x9_y18),
    .I3(x9_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111010000111)
) lut_13_14 (
    .O(x13_y14),
    .I0(1'b0),
    .I1(x10_y13),
    .I2(1'b0),
    .I3(x10_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111100001100)
) lut_14_14 (
    .O(x14_y14),
    .I0(x11_y19),
    .I1(1'b0),
    .I2(x12_y9),
    .I3(x11_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011110101001)
) lut_15_14 (
    .O(x15_y14),
    .I0(1'b0),
    .I1(x13_y12),
    .I2(x12_y12),
    .I3(x13_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011011010111)
) lut_16_14 (
    .O(x16_y14),
    .I0(x14_y12),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x14_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110011010001)
) lut_17_14 (
    .O(x17_y14),
    .I0(x14_y15),
    .I1(x15_y19),
    .I2(x14_y11),
    .I3(x15_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010000110101)
) lut_18_14 (
    .O(x18_y14),
    .I0(1'b0),
    .I1(x16_y13),
    .I2(x15_y14),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100001110101)
) lut_19_14 (
    .O(x19_y14),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001110101000)
) lut_20_14 (
    .O(x20_y14),
    .I0(x18_y19),
    .I1(1'b0),
    .I2(x18_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010110101000)
) lut_21_14 (
    .O(x21_y14),
    .I0(x18_y17),
    .I1(1'b0),
    .I2(x18_y11),
    .I3(x19_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111000000000)
) lut_22_14 (
    .O(x22_y14),
    .I0(1'b0),
    .I1(x20_y10),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110110001111)
) lut_23_14 (
    .O(x23_y14),
    .I0(x20_y13),
    .I1(x21_y15),
    .I2(x21_y9),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101110110000)
) lut_24_14 (
    .O(x24_y14),
    .I0(x22_y19),
    .I1(x22_y10),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111111101110)
) lut_25_14 (
    .O(x25_y14),
    .I0(1'b0),
    .I1(x23_y11),
    .I2(x22_y15),
    .I3(x23_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101001101001)
) lut_26_14 (
    .O(x26_y14),
    .I0(x24_y12),
    .I1(x24_y15),
    .I2(x24_y16),
    .I3(x24_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001000001100)
) lut_27_14 (
    .O(x27_y14),
    .I0(x25_y19),
    .I1(1'b0),
    .I2(x24_y10),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110001110001)
) lut_28_14 (
    .O(x28_y14),
    .I0(x26_y9),
    .I1(x25_y14),
    .I2(1'b0),
    .I3(x26_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110011100011)
) lut_29_14 (
    .O(x29_y14),
    .I0(x27_y9),
    .I1(x26_y12),
    .I2(1'b0),
    .I3(x27_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101001001010)
) lut_30_14 (
    .O(x30_y14),
    .I0(x28_y12),
    .I1(x28_y14),
    .I2(x27_y13),
    .I3(x28_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010001001101)
) lut_31_14 (
    .O(x31_y14),
    .I0(1'b0),
    .I1(x29_y15),
    .I2(x29_y13),
    .I3(x29_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000010101110)
) lut_32_14 (
    .O(x32_y14),
    .I0(x29_y9),
    .I1(x29_y15),
    .I2(x30_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010111110010)
) lut_33_14 (
    .O(x33_y14),
    .I0(x31_y14),
    .I1(x30_y9),
    .I2(x30_y16),
    .I3(x30_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001110001111)
) lut_34_14 (
    .O(x34_y14),
    .I0(x31_y16),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x31_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111000011101)
) lut_35_14 (
    .O(x35_y14),
    .I0(1'b0),
    .I1(x32_y16),
    .I2(x32_y14),
    .I3(x32_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001110011011)
) lut_36_14 (
    .O(x36_y14),
    .I0(x33_y14),
    .I1(x34_y13),
    .I2(x33_y9),
    .I3(x34_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010110000010)
) lut_37_14 (
    .O(x37_y14),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x34_y13),
    .I3(x35_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110100010111)
) lut_38_14 (
    .O(x38_y14),
    .I0(x35_y16),
    .I1(x35_y14),
    .I2(x35_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010100100000)
) lut_39_14 (
    .O(x39_y14),
    .I0(x37_y17),
    .I1(1'b0),
    .I2(x36_y16),
    .I3(x36_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001000011010)
) lut_40_14 (
    .O(x40_y14),
    .I0(x38_y17),
    .I1(x38_y9),
    .I2(1'b0),
    .I3(x37_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001110100001)
) lut_41_14 (
    .O(x41_y14),
    .I0(x39_y13),
    .I1(x38_y9),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001011011100)
) lut_42_14 (
    .O(x42_y14),
    .I0(1'b0),
    .I1(x40_y10),
    .I2(x40_y10),
    .I3(x40_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000100111101)
) lut_43_14 (
    .O(x43_y14),
    .I0(x41_y16),
    .I1(x41_y15),
    .I2(x40_y19),
    .I3(x40_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010110101011)
) lut_44_14 (
    .O(x44_y14),
    .I0(x42_y11),
    .I1(x41_y14),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011000100011)
) lut_45_14 (
    .O(x45_y14),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x43_y13),
    .I3(x43_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011111111001)
) lut_46_14 (
    .O(x46_y14),
    .I0(1'b0),
    .I1(x43_y16),
    .I2(1'b0),
    .I3(x43_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000100000111)
) lut_47_14 (
    .O(x47_y14),
    .I0(1'b0),
    .I1(x44_y16),
    .I2(x44_y11),
    .I3(x45_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111101001000)
) lut_48_14 (
    .O(x48_y14),
    .I0(x46_y9),
    .I1(x46_y12),
    .I2(x45_y10),
    .I3(x46_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100000101101)
) lut_49_14 (
    .O(x49_y14),
    .I0(1'b0),
    .I1(x46_y13),
    .I2(1'b0),
    .I3(x47_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010100010000)
) lut_50_14 (
    .O(x50_y14),
    .I0(x48_y11),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x47_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101000100001)
) lut_51_14 (
    .O(x51_y14),
    .I0(x49_y10),
    .I1(1'b0),
    .I2(x48_y13),
    .I3(x48_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001101011110)
) lut_52_14 (
    .O(x52_y14),
    .I0(1'b0),
    .I1(x49_y9),
    .I2(x49_y11),
    .I3(x49_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111010110101)
) lut_53_14 (
    .O(x53_y14),
    .I0(x51_y15),
    .I1(x51_y9),
    .I2(x51_y16),
    .I3(x51_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101100000110)
) lut_54_14 (
    .O(x54_y14),
    .I0(x51_y10),
    .I1(1'b0),
    .I2(x52_y13),
    .I3(x51_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100111010100)
) lut_55_14 (
    .O(x55_y14),
    .I0(x52_y19),
    .I1(x52_y15),
    .I2(x52_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110111000111)
) lut_56_14 (
    .O(x56_y14),
    .I0(x54_y14),
    .I1(x53_y12),
    .I2(x54_y18),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100011010001)
) lut_57_14 (
    .O(x57_y14),
    .I0(x54_y10),
    .I1(x54_y18),
    .I2(x54_y18),
    .I3(x55_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111110011110)
) lut_58_14 (
    .O(x58_y14),
    .I0(x56_y16),
    .I1(x56_y13),
    .I2(x56_y19),
    .I3(x55_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001011110111)
) lut_59_14 (
    .O(x59_y14),
    .I0(x56_y19),
    .I1(x57_y10),
    .I2(x57_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001100100000)
) lut_60_14 (
    .O(x60_y14),
    .I0(x58_y18),
    .I1(x58_y19),
    .I2(1'b0),
    .I3(x57_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010111001100)
) lut_61_14 (
    .O(x61_y14),
    .I0(x59_y15),
    .I1(x58_y13),
    .I2(x59_y17),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000000100110)
) lut_62_14 (
    .O(x62_y14),
    .I0(x60_y16),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x59_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100001000111)
) lut_0_15 (
    .O(x0_y15),
    .I0(in4),
    .I1(in2),
    .I2(in6),
    .I3(in9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101001100111)
) lut_1_15 (
    .O(x1_y15),
    .I0(in3),
    .I1(in0),
    .I2(in1),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100001000101)
) lut_2_15 (
    .O(x2_y15),
    .I0(in5),
    .I1(in7),
    .I2(1'b0),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100001000111)
) lut_3_15 (
    .O(x3_y15),
    .I0(1'b0),
    .I1(x1_y12),
    .I2(in0),
    .I3(x1_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011100110100)
) lut_4_15 (
    .O(x4_y15),
    .I0(x1_y10),
    .I1(x2_y12),
    .I2(x1_y12),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001100000100)
) lut_5_15 (
    .O(x5_y15),
    .I0(x2_y15),
    .I1(x2_y17),
    .I2(x3_y10),
    .I3(x3_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111100000111)
) lut_6_15 (
    .O(x6_y15),
    .I0(x3_y15),
    .I1(x3_y14),
    .I2(x4_y11),
    .I3(x3_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010100011110)
) lut_7_15 (
    .O(x7_y15),
    .I0(1'b0),
    .I1(x5_y17),
    .I2(x5_y20),
    .I3(x4_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000011110000)
) lut_8_15 (
    .O(x8_y15),
    .I0(1'b0),
    .I1(x6_y11),
    .I2(x6_y11),
    .I3(x6_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000110010110)
) lut_9_15 (
    .O(x9_y15),
    .I0(x6_y16),
    .I1(x6_y20),
    .I2(x6_y11),
    .I3(x6_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101110010110)
) lut_10_15 (
    .O(x10_y15),
    .I0(x8_y18),
    .I1(x7_y19),
    .I2(x8_y12),
    .I3(x7_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011110101000)
) lut_11_15 (
    .O(x11_y15),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x8_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111110111111)
) lut_12_15 (
    .O(x12_y15),
    .I0(x10_y18),
    .I1(x9_y17),
    .I2(x9_y19),
    .I3(x10_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010001011011)
) lut_13_15 (
    .O(x13_y15),
    .I0(1'b0),
    .I1(x11_y10),
    .I2(x11_y17),
    .I3(x10_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110000110101)
) lut_14_15 (
    .O(x14_y15),
    .I0(x11_y18),
    .I1(x12_y11),
    .I2(x11_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011011011011)
) lut_15_15 (
    .O(x15_y15),
    .I0(1'b0),
    .I1(x12_y14),
    .I2(x13_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011100110111)
) lut_16_15 (
    .O(x16_y15),
    .I0(x14_y18),
    .I1(1'b0),
    .I2(x14_y14),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110001110011)
) lut_17_15 (
    .O(x17_y15),
    .I0(1'b0),
    .I1(x15_y18),
    .I2(x15_y13),
    .I3(x14_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101101101011)
) lut_18_15 (
    .O(x18_y15),
    .I0(x16_y11),
    .I1(x16_y10),
    .I2(x15_y12),
    .I3(x16_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001011010111)
) lut_19_15 (
    .O(x19_y15),
    .I0(x17_y18),
    .I1(x16_y18),
    .I2(x16_y20),
    .I3(x17_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011000000011)
) lut_20_15 (
    .O(x20_y15),
    .I0(x17_y12),
    .I1(x17_y13),
    .I2(x17_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111100101000)
) lut_21_15 (
    .O(x21_y15),
    .I0(x18_y14),
    .I1(x19_y13),
    .I2(x18_y15),
    .I3(x18_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010010000000)
) lut_22_15 (
    .O(x22_y15),
    .I0(1'b0),
    .I1(x20_y18),
    .I2(x20_y13),
    .I3(x20_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000000001010)
) lut_23_15 (
    .O(x23_y15),
    .I0(x20_y19),
    .I1(x20_y14),
    .I2(x20_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111011010111)
) lut_24_15 (
    .O(x24_y15),
    .I0(1'b0),
    .I1(x21_y14),
    .I2(1'b0),
    .I3(x22_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010010001110)
) lut_25_15 (
    .O(x25_y15),
    .I0(x22_y16),
    .I1(x23_y20),
    .I2(x23_y20),
    .I3(x22_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000110001110)
) lut_26_15 (
    .O(x26_y15),
    .I0(1'b0),
    .I1(x24_y11),
    .I2(x24_y19),
    .I3(x24_y10)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101001110111)
) lut_27_15 (
    .O(x27_y15),
    .I0(x25_y16),
    .I1(x25_y10),
    .I2(x25_y16),
    .I3(x24_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100011011001)
) lut_28_15 (
    .O(x28_y15),
    .I0(x25_y14),
    .I1(x25_y13),
    .I2(x26_y19),
    .I3(x25_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011100011010)
) lut_29_15 (
    .O(x29_y15),
    .I0(x27_y19),
    .I1(x26_y11),
    .I2(1'b0),
    .I3(x26_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011010011110)
) lut_30_15 (
    .O(x30_y15),
    .I0(x27_y11),
    .I1(x28_y11),
    .I2(x28_y20),
    .I3(x27_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101001101111)
) lut_31_15 (
    .O(x31_y15),
    .I0(x29_y17),
    .I1(1'b0),
    .I2(x29_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001001110110)
) lut_32_15 (
    .O(x32_y15),
    .I0(x29_y15),
    .I1(x29_y14),
    .I2(x29_y14),
    .I3(x30_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111100010001)
) lut_33_15 (
    .O(x33_y15),
    .I0(x31_y12),
    .I1(x31_y11),
    .I2(1'b0),
    .I3(x30_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110000111000)
) lut_34_15 (
    .O(x34_y15),
    .I0(1'b0),
    .I1(x32_y16),
    .I2(x32_y13),
    .I3(x32_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010100111111)
) lut_35_15 (
    .O(x35_y15),
    .I0(x32_y14),
    .I1(x32_y14),
    .I2(x32_y15),
    .I3(x32_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000101111101)
) lut_36_15 (
    .O(x36_y15),
    .I0(1'b0),
    .I1(x33_y17),
    .I2(x34_y15),
    .I3(x33_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011000000110)
) lut_37_15 (
    .O(x37_y15),
    .I0(1'b0),
    .I1(x35_y16),
    .I2(x34_y16),
    .I3(x34_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101101011110)
) lut_38_15 (
    .O(x38_y15),
    .I0(x36_y18),
    .I1(x36_y19),
    .I2(1'b0),
    .I3(x35_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000010110111)
) lut_39_15 (
    .O(x39_y15),
    .I0(x37_y14),
    .I1(x36_y19),
    .I2(1'b0),
    .I3(x37_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000011101011)
) lut_40_15 (
    .O(x40_y15),
    .I0(x38_y11),
    .I1(x38_y17),
    .I2(1'b0),
    .I3(x38_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111100100110)
) lut_41_15 (
    .O(x41_y15),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x38_y16),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111101010100)
) lut_42_15 (
    .O(x42_y15),
    .I0(x39_y15),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x39_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101110001100)
) lut_43_15 (
    .O(x43_y15),
    .I0(x40_y17),
    .I1(1'b0),
    .I2(x40_y18),
    .I3(x41_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100111101101)
) lut_44_15 (
    .O(x44_y15),
    .I0(x41_y13),
    .I1(x41_y16),
    .I2(1'b0),
    .I3(x42_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000011110110)
) lut_45_15 (
    .O(x45_y15),
    .I0(1'b0),
    .I1(x42_y10),
    .I2(1'b0),
    .I3(x42_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101110010110)
) lut_46_15 (
    .O(x46_y15),
    .I0(x44_y10),
    .I1(x43_y19),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001110110101)
) lut_47_15 (
    .O(x47_y15),
    .I0(x45_y10),
    .I1(x45_y12),
    .I2(1'b0),
    .I3(x44_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011001100000)
) lut_48_15 (
    .O(x48_y15),
    .I0(x46_y14),
    .I1(x45_y15),
    .I2(1'b0),
    .I3(x45_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001110110101)
) lut_49_15 (
    .O(x49_y15),
    .I0(x47_y11),
    .I1(x47_y18),
    .I2(x47_y16),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010100110110)
) lut_50_15 (
    .O(x50_y15),
    .I0(x47_y13),
    .I1(x47_y13),
    .I2(x47_y18),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110000110010)
) lut_51_15 (
    .O(x51_y15),
    .I0(x48_y10),
    .I1(x48_y11),
    .I2(x48_y16),
    .I3(x48_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010010101111)
) lut_52_15 (
    .O(x52_y15),
    .I0(x49_y17),
    .I1(x49_y15),
    .I2(1'b0),
    .I3(x50_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110001100100)
) lut_53_15 (
    .O(x53_y15),
    .I0(x51_y14),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100000011111)
) lut_54_15 (
    .O(x54_y15),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x52_y18),
    .I3(x52_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001110000100)
) lut_55_15 (
    .O(x55_y15),
    .I0(x53_y12),
    .I1(x53_y12),
    .I2(x52_y20),
    .I3(x53_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010100111111)
) lut_56_15 (
    .O(x56_y15),
    .I0(x54_y16),
    .I1(x53_y14),
    .I2(x53_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001000001001)
) lut_57_15 (
    .O(x57_y15),
    .I0(x54_y10),
    .I1(x54_y15),
    .I2(x55_y11),
    .I3(x55_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100010000011)
) lut_58_15 (
    .O(x58_y15),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x56_y18),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011010101011)
) lut_59_15 (
    .O(x59_y15),
    .I0(x56_y17),
    .I1(x56_y12),
    .I2(x56_y17),
    .I3(x56_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100101110001)
) lut_60_15 (
    .O(x60_y15),
    .I0(x57_y14),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x58_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111100011000)
) lut_61_15 (
    .O(x61_y15),
    .I0(x59_y14),
    .I1(x58_y10),
    .I2(x58_y10),
    .I3(x58_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001100010100)
) lut_62_15 (
    .O(x62_y15),
    .I0(x59_y14),
    .I1(x59_y18),
    .I2(1'b0),
    .I3(x59_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100001100111)
) lut_0_16 (
    .O(x0_y16),
    .I0(in1),
    .I1(1'b0),
    .I2(in7),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010001010100)
) lut_1_16 (
    .O(x1_y16),
    .I0(in4),
    .I1(in2),
    .I2(in9),
    .I3(in4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001111000110)
) lut_2_16 (
    .O(x2_y16),
    .I0(in0),
    .I1(in2),
    .I2(in6),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110111000000)
) lut_3_16 (
    .O(x3_y16),
    .I0(1'b0),
    .I1(1'b0),
    .I2(in9),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011101100000)
) lut_4_16 (
    .O(x4_y16),
    .I0(x2_y20),
    .I1(x2_y11),
    .I2(x1_y20),
    .I3(x2_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110111111001)
) lut_5_16 (
    .O(x5_y16),
    .I0(x2_y13),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x3_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100011110001)
) lut_6_16 (
    .O(x6_y16),
    .I0(x3_y21),
    .I1(x4_y11),
    .I2(x3_y17),
    .I3(x3_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100001101010)
) lut_7_16 (
    .O(x7_y16),
    .I0(x4_y17),
    .I1(x4_y21),
    .I2(x5_y12),
    .I3(x5_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000000001010)
) lut_8_16 (
    .O(x8_y16),
    .I0(x6_y12),
    .I1(1'b0),
    .I2(x5_y21),
    .I3(x5_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001111110011)
) lut_9_16 (
    .O(x9_y16),
    .I0(x7_y17),
    .I1(1'b0),
    .I2(x5_y21),
    .I3(x5_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101011010101)
) lut_10_16 (
    .O(x10_y16),
    .I0(x8_y19),
    .I1(1'b0),
    .I2(x8_y14),
    .I3(x8_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010100111110)
) lut_11_16 (
    .O(x11_y16),
    .I0(x9_y16),
    .I1(x9_y17),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111001101101)
) lut_12_16 (
    .O(x12_y16),
    .I0(x9_y17),
    .I1(x10_y21),
    .I2(x10_y16),
    .I3(x10_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001100111110)
) lut_13_16 (
    .O(x13_y16),
    .I0(x10_y19),
    .I1(x11_y19),
    .I2(x10_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011110000011)
) lut_14_16 (
    .O(x14_y16),
    .I0(x12_y16),
    .I1(x11_y13),
    .I2(1'b0),
    .I3(x12_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101100011001)
) lut_15_16 (
    .O(x15_y16),
    .I0(x12_y21),
    .I1(x13_y16),
    .I2(x12_y18),
    .I3(x12_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100010001111)
) lut_16_16 (
    .O(x16_y16),
    .I0(x13_y11),
    .I1(x13_y20),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010001010100)
) lut_17_16 (
    .O(x17_y16),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x15_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011110111111)
) lut_18_16 (
    .O(x18_y16),
    .I0(x15_y20),
    .I1(x16_y11),
    .I2(1'b0),
    .I3(x15_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100001000111)
) lut_19_16 (
    .O(x19_y16),
    .I0(x17_y12),
    .I1(x16_y11),
    .I2(x17_y14),
    .I3(x17_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010101110110)
) lut_20_16 (
    .O(x20_y16),
    .I0(x18_y16),
    .I1(x17_y21),
    .I2(x17_y17),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100000001101)
) lut_21_16 (
    .O(x21_y16),
    .I0(x18_y11),
    .I1(x19_y21),
    .I2(x18_y12),
    .I3(x18_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000111011000)
) lut_22_16 (
    .O(x22_y16),
    .I0(1'b0),
    .I1(x19_y21),
    .I2(x20_y20),
    .I3(x20_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101011101010)
) lut_23_16 (
    .O(x23_y16),
    .I0(x21_y16),
    .I1(1'b0),
    .I2(x21_y18),
    .I3(x20_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100101010101)
) lut_24_16 (
    .O(x24_y16),
    .I0(x21_y11),
    .I1(x22_y21),
    .I2(x22_y18),
    .I3(x22_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100000110000)
) lut_25_16 (
    .O(x25_y16),
    .I0(x22_y17),
    .I1(x22_y14),
    .I2(x22_y20),
    .I3(x22_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110011111101)
) lut_26_16 (
    .O(x26_y16),
    .I0(x24_y16),
    .I1(x23_y14),
    .I2(1'b0),
    .I3(x23_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011100000001)
) lut_27_16 (
    .O(x27_y16),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x25_y13),
    .I3(x24_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101001000011)
) lut_28_16 (
    .O(x28_y16),
    .I0(x26_y21),
    .I1(x26_y14),
    .I2(x26_y18),
    .I3(x26_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110101001111)
) lut_29_16 (
    .O(x29_y16),
    .I0(1'b0),
    .I1(x26_y21),
    .I2(1'b0),
    .I3(x27_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010100111100)
) lut_30_16 (
    .O(x30_y16),
    .I0(1'b0),
    .I1(x27_y11),
    .I2(x27_y12),
    .I3(x27_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000010101101)
) lut_31_16 (
    .O(x31_y16),
    .I0(x28_y16),
    .I1(x29_y14),
    .I2(x29_y16),
    .I3(x28_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000101111011)
) lut_32_16 (
    .O(x32_y16),
    .I0(x30_y19),
    .I1(1'b0),
    .I2(x29_y11),
    .I3(x29_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100001011110)
) lut_33_16 (
    .O(x33_y16),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x30_y19),
    .I3(x30_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001100000000)
) lut_34_16 (
    .O(x34_y16),
    .I0(x32_y16),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x31_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000110001110)
) lut_35_16 (
    .O(x35_y16),
    .I0(x33_y20),
    .I1(x33_y18),
    .I2(x33_y11),
    .I3(x33_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011101000101)
) lut_36_16 (
    .O(x36_y16),
    .I0(x34_y11),
    .I1(x34_y16),
    .I2(x33_y21),
    .I3(x33_y11)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111011111010)
) lut_37_16 (
    .O(x37_y16),
    .I0(x35_y11),
    .I1(x34_y14),
    .I2(1'b0),
    .I3(x35_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001001000010)
) lut_38_16 (
    .O(x38_y16),
    .I0(x36_y21),
    .I1(x35_y15),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011100101111)
) lut_39_16 (
    .O(x39_y16),
    .I0(x37_y18),
    .I1(x36_y20),
    .I2(x37_y18),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000101111000)
) lut_40_16 (
    .O(x40_y16),
    .I0(x37_y20),
    .I1(x37_y16),
    .I2(1'b0),
    .I3(x37_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001110001110)
) lut_41_16 (
    .O(x41_y16),
    .I0(x38_y14),
    .I1(x39_y13),
    .I2(1'b0),
    .I3(x39_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010001001000)
) lut_42_16 (
    .O(x42_y16),
    .I0(x39_y19),
    .I1(1'b0),
    .I2(x40_y16),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010001100000)
) lut_43_16 (
    .O(x43_y16),
    .I0(x41_y11),
    .I1(x40_y18),
    .I2(x40_y14),
    .I3(x41_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001101100111)
) lut_44_16 (
    .O(x44_y16),
    .I0(x42_y21),
    .I1(x42_y20),
    .I2(x42_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111110001111)
) lut_45_16 (
    .O(x45_y16),
    .I0(x42_y15),
    .I1(1'b0),
    .I2(x42_y13),
    .I3(x42_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111010001000)
) lut_46_16 (
    .O(x46_y16),
    .I0(x43_y20),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110010100000)
) lut_47_16 (
    .O(x47_y16),
    .I0(x45_y20),
    .I1(x45_y15),
    .I2(1'b0),
    .I3(x44_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001000010110)
) lut_48_16 (
    .O(x48_y16),
    .I0(x46_y14),
    .I1(x46_y19),
    .I2(x46_y20),
    .I3(x46_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011100110011)
) lut_49_16 (
    .O(x49_y16),
    .I0(x47_y17),
    .I1(x47_y19),
    .I2(1'b0),
    .I3(x46_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100000001101)
) lut_50_16 (
    .O(x50_y16),
    .I0(x47_y16),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x47_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111101001111)
) lut_51_16 (
    .O(x51_y16),
    .I0(1'b0),
    .I1(x49_y12),
    .I2(1'b0),
    .I3(x49_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000001100111)
) lut_52_16 (
    .O(x52_y16),
    .I0(x50_y15),
    .I1(x49_y11),
    .I2(x49_y16),
    .I3(x49_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101011110010)
) lut_53_16 (
    .O(x53_y16),
    .I0(x51_y14),
    .I1(1'b0),
    .I2(x51_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110110110111)
) lut_54_16 (
    .O(x54_y16),
    .I0(x51_y11),
    .I1(x51_y21),
    .I2(x52_y21),
    .I3(x52_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111111111001)
) lut_55_16 (
    .O(x55_y16),
    .I0(x52_y14),
    .I1(x52_y16),
    .I2(x52_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001011001001)
) lut_56_16 (
    .O(x56_y16),
    .I0(x54_y18),
    .I1(1'b0),
    .I2(x53_y11),
    .I3(x54_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110111100110)
) lut_57_16 (
    .O(x57_y16),
    .I0(x54_y19),
    .I1(x54_y14),
    .I2(x54_y14),
    .I3(x54_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011110000010)
) lut_58_16 (
    .O(x58_y16),
    .I0(x56_y17),
    .I1(1'b0),
    .I2(x56_y14),
    .I3(x55_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101000000001)
) lut_59_16 (
    .O(x59_y16),
    .I0(x57_y13),
    .I1(x57_y21),
    .I2(1'b0),
    .I3(x57_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111101000011)
) lut_60_16 (
    .O(x60_y16),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x57_y20),
    .I3(x58_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111110000001)
) lut_61_16 (
    .O(x61_y16),
    .I0(x59_y21),
    .I1(1'b0),
    .I2(x59_y18),
    .I3(x59_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010000110010)
) lut_62_16 (
    .O(x62_y16),
    .I0(x60_y11),
    .I1(x60_y16),
    .I2(x59_y15),
    .I3(x59_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000111010110)
) lut_0_17 (
    .O(x0_y17),
    .I0(in9),
    .I1(in5),
    .I2(1'b0),
    .I3(in4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011000011000)
) lut_1_17 (
    .O(x1_y17),
    .I0(1'b0),
    .I1(in8),
    .I2(in8),
    .I3(in4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111000101110)
) lut_2_17 (
    .O(x2_y17),
    .I0(in3),
    .I1(1'b0),
    .I2(1'b0),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011111011110)
) lut_3_17 (
    .O(x3_y17),
    .I0(in8),
    .I1(1'b0),
    .I2(in1),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111011110100)
) lut_4_17 (
    .O(x4_y17),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x1_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000001101101)
) lut_5_17 (
    .O(x5_y17),
    .I0(x2_y15),
    .I1(x3_y13),
    .I2(1'b0),
    .I3(x3_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010100110101)
) lut_6_17 (
    .O(x6_y17),
    .I0(x3_y16),
    .I1(x3_y19),
    .I2(x4_y14),
    .I3(x4_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100101001001)
) lut_7_17 (
    .O(x7_y17),
    .I0(x4_y16),
    .I1(x4_y19),
    .I2(x5_y21),
    .I3(x5_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001110110101)
) lut_8_17 (
    .O(x8_y17),
    .I0(x6_y17),
    .I1(x5_y21),
    .I2(x6_y16),
    .I3(x5_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000000000010)
) lut_9_17 (
    .O(x9_y17),
    .I0(x6_y19),
    .I1(x7_y20),
    .I2(x6_y16),
    .I3(x5_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110010100000)
) lut_10_17 (
    .O(x10_y17),
    .I0(x7_y16),
    .I1(x7_y20),
    .I2(x7_y14),
    .I3(x7_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001100101000)
) lut_11_17 (
    .O(x11_y17),
    .I0(x8_y18),
    .I1(x9_y22),
    .I2(x8_y19),
    .I3(x9_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001000010110)
) lut_12_17 (
    .O(x12_y17),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x9_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011011110111)
) lut_13_17 (
    .O(x13_y17),
    .I0(x11_y18),
    .I1(x10_y13),
    .I2(x11_y15),
    .I3(x11_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000000100001)
) lut_14_17 (
    .O(x14_y17),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x12_y21),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101010010000)
) lut_15_17 (
    .O(x15_y17),
    .I0(x12_y22),
    .I1(x12_y17),
    .I2(1'b0),
    .I3(x12_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101001100011)
) lut_16_17 (
    .O(x16_y17),
    .I0(1'b0),
    .I1(x13_y16),
    .I2(x14_y17),
    .I3(x14_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101010111110)
) lut_17_17 (
    .O(x17_y17),
    .I0(x15_y20),
    .I1(1'b0),
    .I2(x15_y20),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000111001100)
) lut_18_17 (
    .O(x18_y17),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x16_y17),
    .I3(x15_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101110011100)
) lut_19_17 (
    .O(x19_y17),
    .I0(x17_y22),
    .I1(1'b0),
    .I2(x17_y15),
    .I3(x17_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110100100000)
) lut_20_17 (
    .O(x20_y17),
    .I0(1'b0),
    .I1(x17_y22),
    .I2(x17_y17),
    .I3(x17_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111010011010)
) lut_21_17 (
    .O(x21_y17),
    .I0(x18_y18),
    .I1(x19_y18),
    .I2(x18_y14),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000011011010)
) lut_22_17 (
    .O(x22_y17),
    .I0(x20_y20),
    .I1(1'b0),
    .I2(x20_y13),
    .I3(x20_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001001000000)
) lut_23_17 (
    .O(x23_y17),
    .I0(x20_y17),
    .I1(x20_y13),
    .I2(x20_y19),
    .I3(x20_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010111110011)
) lut_24_17 (
    .O(x24_y17),
    .I0(x22_y13),
    .I1(x22_y22),
    .I2(x22_y18),
    .I3(x21_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100101011100)
) lut_25_17 (
    .O(x25_y17),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x23_y21),
    .I3(x22_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110010101100)
) lut_26_17 (
    .O(x26_y17),
    .I0(x24_y20),
    .I1(x23_y18),
    .I2(x23_y19),
    .I3(x24_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010111010110)
) lut_27_17 (
    .O(x27_y17),
    .I0(x25_y15),
    .I1(x24_y16),
    .I2(x24_y13),
    .I3(x25_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111011011010)
) lut_28_17 (
    .O(x28_y17),
    .I0(x26_y18),
    .I1(1'b0),
    .I2(x26_y16),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011110010011)
) lut_29_17 (
    .O(x29_y17),
    .I0(x26_y21),
    .I1(x26_y18),
    .I2(1'b0),
    .I3(x27_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000001111101)
) lut_30_17 (
    .O(x30_y17),
    .I0(1'b0),
    .I1(x27_y17),
    .I2(x27_y22),
    .I3(x27_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111101100111)
) lut_31_17 (
    .O(x31_y17),
    .I0(1'b0),
    .I1(x28_y14),
    .I2(x28_y20),
    .I3(x29_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100100001100)
) lut_32_17 (
    .O(x32_y17),
    .I0(1'b0),
    .I1(x29_y16),
    .I2(1'b0),
    .I3(x30_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001001110100)
) lut_33_17 (
    .O(x33_y17),
    .I0(x30_y21),
    .I1(x30_y17),
    .I2(x31_y19),
    .I3(x30_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010101111111)
) lut_34_17 (
    .O(x34_y17),
    .I0(x32_y22),
    .I1(x32_y19),
    .I2(x31_y21),
    .I3(x31_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011100101111)
) lut_35_17 (
    .O(x35_y17),
    .I0(x33_y22),
    .I1(x32_y13),
    .I2(x32_y18),
    .I3(x32_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110011000010)
) lut_36_17 (
    .O(x36_y17),
    .I0(x33_y21),
    .I1(1'b0),
    .I2(x34_y18),
    .I3(x33_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000111110101)
) lut_37_17 (
    .O(x37_y17),
    .I0(x34_y12),
    .I1(x34_y19),
    .I2(x34_y12),
    .I3(x34_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011100000110)
) lut_38_17 (
    .O(x38_y17),
    .I0(1'b0),
    .I1(x36_y14),
    .I2(1'b0),
    .I3(x35_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110011011011)
) lut_39_17 (
    .O(x39_y17),
    .I0(1'b0),
    .I1(x37_y14),
    .I2(x36_y19),
    .I3(x37_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110000010110)
) lut_40_17 (
    .O(x40_y17),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x38_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000011100010)
) lut_41_17 (
    .O(x41_y17),
    .I0(x39_y17),
    .I1(x39_y14),
    .I2(1'b0),
    .I3(x38_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011011110100)
) lut_42_17 (
    .O(x42_y17),
    .I0(x39_y16),
    .I1(x39_y18),
    .I2(1'b0),
    .I3(x40_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111001011111)
) lut_43_17 (
    .O(x43_y17),
    .I0(x40_y15),
    .I1(1'b0),
    .I2(x41_y17),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000110000111)
) lut_44_17 (
    .O(x44_y17),
    .I0(x41_y17),
    .I1(1'b0),
    .I2(x42_y19),
    .I3(x41_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010101100011)
) lut_45_17 (
    .O(x45_y17),
    .I0(1'b0),
    .I1(x42_y18),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010101001101)
) lut_46_17 (
    .O(x46_y17),
    .I0(x44_y18),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000100101011)
) lut_47_17 (
    .O(x47_y17),
    .I0(x44_y19),
    .I1(x44_y14),
    .I2(1'b0),
    .I3(x45_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011101001001)
) lut_48_17 (
    .O(x48_y17),
    .I0(x46_y14),
    .I1(x45_y17),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111100111011)
) lut_49_17 (
    .O(x49_y17),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x46_y15),
    .I3(x46_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100100111001)
) lut_50_17 (
    .O(x50_y17),
    .I0(1'b0),
    .I1(x48_y21),
    .I2(1'b0),
    .I3(x48_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110100111101)
) lut_51_17 (
    .O(x51_y17),
    .I0(x49_y19),
    .I1(x48_y16),
    .I2(x49_y12),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010100111100)
) lut_52_17 (
    .O(x52_y17),
    .I0(1'b0),
    .I1(x49_y12),
    .I2(1'b0),
    .I3(x49_y12)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011010011101)
) lut_53_17 (
    .O(x53_y17),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x51_y13),
    .I3(x51_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100111101001)
) lut_54_17 (
    .O(x54_y17),
    .I0(x51_y12),
    .I1(x52_y21),
    .I2(1'b0),
    .I3(x51_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000100110001)
) lut_55_17 (
    .O(x55_y17),
    .I0(x53_y13),
    .I1(x52_y20),
    .I2(x53_y15),
    .I3(x52_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011101011111)
) lut_56_17 (
    .O(x56_y17),
    .I0(x53_y14),
    .I1(1'b0),
    .I2(x54_y17),
    .I3(x53_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010100100110)
) lut_57_17 (
    .O(x57_y17),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x54_y14),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110011011110)
) lut_58_17 (
    .O(x58_y17),
    .I0(x56_y19),
    .I1(x55_y19),
    .I2(1'b0),
    .I3(x55_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001101010111)
) lut_59_17 (
    .O(x59_y17),
    .I0(x57_y21),
    .I1(x56_y20),
    .I2(x57_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001000010011)
) lut_60_17 (
    .O(x60_y17),
    .I0(x58_y14),
    .I1(1'b0),
    .I2(x58_y18),
    .I3(x57_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011100000011)
) lut_61_17 (
    .O(x61_y17),
    .I0(x59_y17),
    .I1(x59_y21),
    .I2(x58_y13),
    .I3(x59_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100110100100)
) lut_62_17 (
    .O(x62_y17),
    .I0(x59_y19),
    .I1(1'b0),
    .I2(x60_y19),
    .I3(x60_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011010100111)
) lut_0_18 (
    .O(x0_y18),
    .I0(1'b0),
    .I1(in1),
    .I2(in8),
    .I3(in4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100110100001)
) lut_1_18 (
    .O(x1_y18),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111001000011)
) lut_2_18 (
    .O(x2_y18),
    .I0(in5),
    .I1(in7),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001000000000)
) lut_3_18 (
    .O(x3_y18),
    .I0(1'b0),
    .I1(in8),
    .I2(in5),
    .I3(x1_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100100111110)
) lut_4_18 (
    .O(x4_y18),
    .I0(x1_y17),
    .I1(x1_y15),
    .I2(x1_y18),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010000000001)
) lut_5_18 (
    .O(x5_y18),
    .I0(x3_y19),
    .I1(1'b0),
    .I2(x2_y19),
    .I3(x2_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111011101000)
) lut_6_18 (
    .O(x6_y18),
    .I0(x4_y17),
    .I1(x4_y20),
    .I2(x3_y14),
    .I3(x3_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010111011011)
) lut_7_18 (
    .O(x7_y18),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x5_y23),
    .I3(x5_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101001111010)
) lut_8_18 (
    .O(x8_y18),
    .I0(1'b0),
    .I1(x5_y13),
    .I2(x6_y23),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111011001001)
) lut_9_18 (
    .O(x9_y18),
    .I0(x6_y20),
    .I1(x7_y15),
    .I2(x6_y23),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110100000110)
) lut_10_18 (
    .O(x10_y18),
    .I0(x8_y21),
    .I1(x8_y15),
    .I2(x8_y14),
    .I3(x8_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110011011111)
) lut_11_18 (
    .O(x11_y18),
    .I0(x8_y15),
    .I1(x9_y17),
    .I2(x9_y16),
    .I3(x8_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000100011000)
) lut_12_18 (
    .O(x12_y18),
    .I0(x10_y16),
    .I1(x9_y14),
    .I2(x9_y21),
    .I3(x10_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111101010001)
) lut_13_18 (
    .O(x13_y18),
    .I0(x10_y17),
    .I1(1'b0),
    .I2(x10_y18),
    .I3(x11_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011100111010)
) lut_14_18 (
    .O(x14_y18),
    .I0(x12_y20),
    .I1(x11_y18),
    .I2(x11_y17),
    .I3(x11_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000001100000)
) lut_15_18 (
    .O(x15_y18),
    .I0(x12_y19),
    .I1(x13_y21),
    .I2(x13_y21),
    .I3(x12_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000100101010)
) lut_16_18 (
    .O(x16_y18),
    .I0(x13_y23),
    .I1(x14_y16),
    .I2(x13_y21),
    .I3(x14_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000011111000)
) lut_17_18 (
    .O(x17_y18),
    .I0(x14_y23),
    .I1(x14_y22),
    .I2(x15_y23),
    .I3(x15_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000100011101)
) lut_18_18 (
    .O(x18_y18),
    .I0(x15_y23),
    .I1(x16_y13),
    .I2(x15_y20),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001001101010)
) lut_19_18 (
    .O(x19_y18),
    .I0(1'b0),
    .I1(x16_y20),
    .I2(x17_y14),
    .I3(x17_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010011010001)
) lut_20_18 (
    .O(x20_y18),
    .I0(x17_y22),
    .I1(x18_y16),
    .I2(1'b0),
    .I3(x17_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100010100100)
) lut_21_18 (
    .O(x21_y18),
    .I0(x18_y23),
    .I1(x18_y17),
    .I2(x18_y17),
    .I3(x19_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110100111010)
) lut_22_18 (
    .O(x22_y18),
    .I0(1'b0),
    .I1(x19_y13),
    .I2(x19_y15),
    .I3(x19_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010011100101)
) lut_23_18 (
    .O(x23_y18),
    .I0(x20_y16),
    .I1(1'b0),
    .I2(x20_y21),
    .I3(x21_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011001011010)
) lut_24_18 (
    .O(x24_y18),
    .I0(x21_y22),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x21_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111010100101)
) lut_25_18 (
    .O(x25_y18),
    .I0(x23_y19),
    .I1(x22_y22),
    .I2(x22_y20),
    .I3(x22_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110100100110)
) lut_26_18 (
    .O(x26_y18),
    .I0(x24_y16),
    .I1(x23_y17),
    .I2(x24_y23),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011010100100)
) lut_27_18 (
    .O(x27_y18),
    .I0(x24_y13),
    .I1(x24_y17),
    .I2(x24_y17),
    .I3(x25_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110110110001)
) lut_28_18 (
    .O(x28_y18),
    .I0(1'b0),
    .I1(x25_y20),
    .I2(1'b0),
    .I3(x25_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100100110010)
) lut_29_18 (
    .O(x29_y18),
    .I0(x27_y16),
    .I1(x27_y23),
    .I2(x27_y16),
    .I3(x27_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000010000110)
) lut_30_18 (
    .O(x30_y18),
    .I0(x28_y20),
    .I1(x28_y21),
    .I2(x28_y19),
    .I3(x28_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100100000100)
) lut_31_18 (
    .O(x31_y18),
    .I0(x28_y15),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x29_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101100101111)
) lut_32_18 (
    .O(x32_y18),
    .I0(x30_y17),
    .I1(x29_y21),
    .I2(x30_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110111011000)
) lut_33_18 (
    .O(x33_y18),
    .I0(x30_y14),
    .I1(x30_y20),
    .I2(x30_y18),
    .I3(x31_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000100001010)
) lut_34_18 (
    .O(x34_y18),
    .I0(1'b0),
    .I1(x31_y17),
    .I2(x32_y22),
    .I3(x31_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010001101111)
) lut_35_18 (
    .O(x35_y18),
    .I0(x32_y20),
    .I1(1'b0),
    .I2(x33_y14),
    .I3(x32_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000011100010)
) lut_36_18 (
    .O(x36_y18),
    .I0(x33_y18),
    .I1(x34_y19),
    .I2(x33_y20),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111111100011)
) lut_37_18 (
    .O(x37_y18),
    .I0(x34_y13),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011100011001)
) lut_38_18 (
    .O(x38_y18),
    .I0(1'b0),
    .I1(x36_y18),
    .I2(1'b0),
    .I3(x35_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000110100001)
) lut_39_18 (
    .O(x39_y18),
    .I0(x37_y14),
    .I1(x37_y22),
    .I2(x37_y21),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011101100011)
) lut_40_18 (
    .O(x40_y18),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x37_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000001010101)
) lut_41_18 (
    .O(x41_y18),
    .I0(x39_y16),
    .I1(x39_y22),
    .I2(x39_y14),
    .I3(x39_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011011101010)
) lut_42_18 (
    .O(x42_y18),
    .I0(x39_y22),
    .I1(x40_y20),
    .I2(x40_y22),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011100001001)
) lut_43_18 (
    .O(x43_y18),
    .I0(x40_y23),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x40_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001010010010)
) lut_44_18 (
    .O(x44_y18),
    .I0(x41_y16),
    .I1(1'b0),
    .I2(x41_y22),
    .I3(x41_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101000000010)
) lut_45_18 (
    .O(x45_y18),
    .I0(x42_y19),
    .I1(x43_y20),
    .I2(x42_y19),
    .I3(x43_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000111101001)
) lut_46_18 (
    .O(x46_y18),
    .I0(x44_y20),
    .I1(x43_y13),
    .I2(x43_y13),
    .I3(x43_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111001010011)
) lut_47_18 (
    .O(x47_y18),
    .I0(1'b0),
    .I1(x44_y13),
    .I2(x44_y16),
    .I3(x44_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100011111110)
) lut_48_18 (
    .O(x48_y18),
    .I0(x46_y16),
    .I1(x46_y19),
    .I2(1'b0),
    .I3(x45_y13)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011110010101)
) lut_49_18 (
    .O(x49_y18),
    .I0(x46_y23),
    .I1(x46_y23),
    .I2(x47_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111101101100)
) lut_50_18 (
    .O(x50_y18),
    .I0(x48_y17),
    .I1(x47_y23),
    .I2(x47_y18),
    .I3(x47_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011001011010)
) lut_51_18 (
    .O(x51_y18),
    .I0(x48_y13),
    .I1(x49_y17),
    .I2(x48_y19),
    .I3(x48_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001010110111)
) lut_52_18 (
    .O(x52_y18),
    .I0(1'b0),
    .I1(x49_y22),
    .I2(x49_y16),
    .I3(x50_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110001010000)
) lut_53_18 (
    .O(x53_y18),
    .I0(x51_y18),
    .I1(x50_y22),
    .I2(x51_y20),
    .I3(x50_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100001001010)
) lut_54_18 (
    .O(x54_y18),
    .I0(x51_y14),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x51_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011100000000)
) lut_55_18 (
    .O(x55_y18),
    .I0(x53_y22),
    .I1(x52_y17),
    .I2(x52_y22),
    .I3(x53_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000010101010)
) lut_56_18 (
    .O(x56_y18),
    .I0(x53_y14),
    .I1(x54_y13),
    .I2(x53_y14),
    .I3(x53_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100001011001)
) lut_57_18 (
    .O(x57_y18),
    .I0(x55_y15),
    .I1(1'b0),
    .I2(x55_y21),
    .I3(x54_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000010101100)
) lut_58_18 (
    .O(x58_y18),
    .I0(1'b0),
    .I1(x56_y18),
    .I2(x56_y16),
    .I3(x56_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010000100000)
) lut_59_18 (
    .O(x59_y18),
    .I0(x57_y13),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x56_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010010011101)
) lut_60_18 (
    .O(x60_y18),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x58_y23),
    .I3(x57_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101001111101)
) lut_61_18 (
    .O(x61_y18),
    .I0(x58_y15),
    .I1(1'b0),
    .I2(x59_y14),
    .I3(x58_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111000110011)
) lut_62_18 (
    .O(x62_y18),
    .I0(x59_y16),
    .I1(1'b0),
    .I2(x59_y22),
    .I3(x59_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101001100000)
) lut_0_19 (
    .O(x0_y19),
    .I0(in8),
    .I1(in3),
    .I2(in0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011011101100)
) lut_1_19 (
    .O(x1_y19),
    .I0(in8),
    .I1(in9),
    .I2(in1),
    .I3(in4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001011010110)
) lut_2_19 (
    .O(x2_y19),
    .I0(in4),
    .I1(1'b0),
    .I2(in6),
    .I3(in4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010111101111)
) lut_3_19 (
    .O(x3_y19),
    .I0(x1_y16),
    .I1(x1_y14),
    .I2(in6),
    .I3(x1_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000111100011)
) lut_4_19 (
    .O(x4_y19),
    .I0(x2_y18),
    .I1(x2_y14),
    .I2(1'b0),
    .I3(x2_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110111010111)
) lut_5_19 (
    .O(x5_y19),
    .I0(x3_y19),
    .I1(x3_y23),
    .I2(x2_y23),
    .I3(x2_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000011111011)
) lut_6_19 (
    .O(x6_y19),
    .I0(x4_y20),
    .I1(1'b0),
    .I2(x3_y17),
    .I3(x4_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010110001110)
) lut_7_19 (
    .O(x7_y19),
    .I0(x4_y15),
    .I1(x4_y22),
    .I2(x5_y23),
    .I3(x5_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001010111001)
) lut_8_19 (
    .O(x8_y19),
    .I0(x5_y20),
    .I1(x6_y19),
    .I2(1'b0),
    .I3(x6_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101011110101)
) lut_9_19 (
    .O(x9_y19),
    .I0(x6_y19),
    .I1(x6_y24),
    .I2(1'b0),
    .I3(x6_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110011101101)
) lut_10_19 (
    .O(x10_y19),
    .I0(x8_y17),
    .I1(x7_y18),
    .I2(x8_y16),
    .I3(x8_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011011101111)
) lut_11_19 (
    .O(x11_y19),
    .I0(x8_y22),
    .I1(x9_y24),
    .I2(x9_y22),
    .I3(x8_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010110101001)
) lut_12_19 (
    .O(x12_y19),
    .I0(x9_y14),
    .I1(x10_y21),
    .I2(x10_y18),
    .I3(x9_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100100011110)
) lut_13_19 (
    .O(x13_y19),
    .I0(1'b0),
    .I1(x10_y15),
    .I2(x11_y19),
    .I3(x10_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100111101011)
) lut_14_19 (
    .O(x14_y19),
    .I0(x12_y22),
    .I1(x12_y24),
    .I2(x11_y23),
    .I3(x11_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101100000000)
) lut_15_19 (
    .O(x15_y19),
    .I0(x12_y20),
    .I1(x12_y16),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101111000001)
) lut_16_19 (
    .O(x16_y19),
    .I0(1'b0),
    .I1(x14_y20),
    .I2(x13_y18),
    .I3(x13_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001001000100)
) lut_17_19 (
    .O(x17_y19),
    .I0(x15_y17),
    .I1(x14_y19),
    .I2(x14_y21),
    .I3(x14_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100011110000)
) lut_18_19 (
    .O(x18_y19),
    .I0(1'b0),
    .I1(x15_y14),
    .I2(1'b0),
    .I3(x16_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100101000111)
) lut_19_19 (
    .O(x19_y19),
    .I0(x16_y17),
    .I1(x16_y22),
    .I2(x16_y17),
    .I3(x17_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000011000010)
) lut_20_19 (
    .O(x20_y19),
    .I0(x18_y22),
    .I1(x18_y15),
    .I2(1'b0),
    .I3(x18_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011001001111)
) lut_21_19 (
    .O(x21_y19),
    .I0(x19_y15),
    .I1(x19_y24),
    .I2(x18_y24),
    .I3(x19_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000000001100)
) lut_22_19 (
    .O(x22_y19),
    .I0(1'b0),
    .I1(x20_y14),
    .I2(x20_y14),
    .I3(x19_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001000011011)
) lut_23_19 (
    .O(x23_y19),
    .I0(x20_y16),
    .I1(x21_y20),
    .I2(x20_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111110101101)
) lut_24_19 (
    .O(x24_y19),
    .I0(x22_y14),
    .I1(1'b0),
    .I2(x21_y14),
    .I3(x22_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100100100001)
) lut_25_19 (
    .O(x25_y19),
    .I0(x22_y19),
    .I1(x23_y23),
    .I2(x23_y22),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001000001011)
) lut_26_19 (
    .O(x26_y19),
    .I0(1'b0),
    .I1(x24_y20),
    .I2(x24_y24),
    .I3(x24_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100111101101)
) lut_27_19 (
    .O(x27_y19),
    .I0(x24_y24),
    .I1(x25_y24),
    .I2(1'b0),
    .I3(x25_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111101101111)
) lut_28_19 (
    .O(x28_y19),
    .I0(1'b0),
    .I1(x25_y23),
    .I2(x26_y14),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101100110000)
) lut_29_19 (
    .O(x29_y19),
    .I0(x26_y21),
    .I1(x27_y21),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010001110011)
) lut_30_19 (
    .O(x30_y19),
    .I0(x27_y20),
    .I1(x27_y16),
    .I2(x28_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010110001100)
) lut_31_19 (
    .O(x31_y19),
    .I0(x28_y19),
    .I1(x28_y22),
    .I2(x29_y21),
    .I3(x28_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001000000100)
) lut_32_19 (
    .O(x32_y19),
    .I0(x30_y19),
    .I1(x30_y16),
    .I2(x29_y24),
    .I3(x29_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011111001101)
) lut_33_19 (
    .O(x33_y19),
    .I0(1'b0),
    .I1(x31_y18),
    .I2(x30_y23),
    .I3(x30_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111011001100)
) lut_34_19 (
    .O(x34_y19),
    .I0(1'b0),
    .I1(x31_y17),
    .I2(x32_y17),
    .I3(x32_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111111110110)
) lut_35_19 (
    .O(x35_y19),
    .I0(x32_y17),
    .I1(x33_y17),
    .I2(x32_y19),
    .I3(x33_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100110100000)
) lut_36_19 (
    .O(x36_y19),
    .I0(x33_y23),
    .I1(1'b0),
    .I2(x33_y17),
    .I3(x34_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111100111100)
) lut_37_19 (
    .O(x37_y19),
    .I0(x34_y14),
    .I1(1'b0),
    .I2(x35_y20),
    .I3(x35_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100101001101)
) lut_38_19 (
    .O(x38_y19),
    .I0(x36_y16),
    .I1(1'b0),
    .I2(x36_y24),
    .I3(x35_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011000101000)
) lut_39_19 (
    .O(x39_y19),
    .I0(x37_y20),
    .I1(x36_y15),
    .I2(x37_y16),
    .I3(x37_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100000111011)
) lut_40_19 (
    .O(x40_y19),
    .I0(1'b0),
    .I1(x38_y14),
    .I2(x38_y24),
    .I3(x37_y14)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011100111100)
) lut_41_19 (
    .O(x41_y19),
    .I0(x39_y16),
    .I1(x39_y23),
    .I2(x39_y24),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010000100110)
) lut_42_19 (
    .O(x42_y19),
    .I0(1'b0),
    .I1(x40_y19),
    .I2(x40_y20),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101110000100)
) lut_43_19 (
    .O(x43_y19),
    .I0(x40_y18),
    .I1(1'b0),
    .I2(x41_y20),
    .I3(x40_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101111101011)
) lut_44_19 (
    .O(x44_y19),
    .I0(x42_y24),
    .I1(x41_y18),
    .I2(x41_y18),
    .I3(x41_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100110100101)
) lut_45_19 (
    .O(x45_y19),
    .I0(x42_y22),
    .I1(x43_y20),
    .I2(x42_y23),
    .I3(x42_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010001011101)
) lut_46_19 (
    .O(x46_y19),
    .I0(x44_y15),
    .I1(x43_y17),
    .I2(x43_y22),
    .I3(x44_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110001110010)
) lut_47_19 (
    .O(x47_y19),
    .I0(x45_y23),
    .I1(x44_y23),
    .I2(x44_y22),
    .I3(x44_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100100000000)
) lut_48_19 (
    .O(x48_y19),
    .I0(x45_y18),
    .I1(x46_y19),
    .I2(x45_y24),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011001011001)
) lut_49_19 (
    .O(x49_y19),
    .I0(x47_y18),
    .I1(x47_y17),
    .I2(x46_y16),
    .I3(x47_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101100001000)
) lut_50_19 (
    .O(x50_y19),
    .I0(x48_y18),
    .I1(x48_y22),
    .I2(x48_y18),
    .I3(x48_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100000101010)
) lut_51_19 (
    .O(x51_y19),
    .I0(x48_y23),
    .I1(x48_y19),
    .I2(x49_y20),
    .I3(x49_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010001001010)
) lut_52_19 (
    .O(x52_y19),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100010011111)
) lut_53_19 (
    .O(x53_y19),
    .I0(x51_y14),
    .I1(x51_y21),
    .I2(x51_y16),
    .I3(x51_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000010011000)
) lut_54_19 (
    .O(x54_y19),
    .I0(x51_y23),
    .I1(x52_y18),
    .I2(1'b0),
    .I3(x52_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010100001001)
) lut_55_19 (
    .O(x55_y19),
    .I0(x53_y23),
    .I1(x53_y22),
    .I2(x52_y20),
    .I3(x52_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111110000101)
) lut_56_19 (
    .O(x56_y19),
    .I0(1'b0),
    .I1(x53_y18),
    .I2(x53_y21),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101010101100)
) lut_57_19 (
    .O(x57_y19),
    .I0(x55_y23),
    .I1(x54_y22),
    .I2(1'b0),
    .I3(x54_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001110000110)
) lut_58_19 (
    .O(x58_y19),
    .I0(x55_y20),
    .I1(x56_y20),
    .I2(1'b0),
    .I3(x56_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101000010110)
) lut_59_19 (
    .O(x59_y19),
    .I0(x56_y19),
    .I1(1'b0),
    .I2(x57_y19),
    .I3(x57_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100001000011)
) lut_60_19 (
    .O(x60_y19),
    .I0(1'b0),
    .I1(x57_y17),
    .I2(x57_y20),
    .I3(x57_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111110111001)
) lut_61_19 (
    .O(x61_y19),
    .I0(x59_y22),
    .I1(x58_y15),
    .I2(x59_y18),
    .I3(x59_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101101110111)
) lut_62_19 (
    .O(x62_y19),
    .I0(x59_y20),
    .I1(x59_y23),
    .I2(1'b0),
    .I3(x60_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110010110000)
) lut_0_20 (
    .O(x0_y20),
    .I0(1'b0),
    .I1(in7),
    .I2(1'b0),
    .I3(in3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000110010011)
) lut_1_20 (
    .O(x1_y20),
    .I0(in9),
    .I1(in9),
    .I2(in5),
    .I3(in4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111110110101)
) lut_2_20 (
    .O(x2_y20),
    .I0(in5),
    .I1(in5),
    .I2(1'b0),
    .I3(in1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011010111101)
) lut_3_20 (
    .O(x3_y20),
    .I0(x1_y23),
    .I1(1'b0),
    .I2(in5),
    .I3(in1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111110010000)
) lut_4_20 (
    .O(x4_y20),
    .I0(x2_y25),
    .I1(x1_y21),
    .I2(1'b0),
    .I3(x1_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101110110001)
) lut_5_20 (
    .O(x5_y20),
    .I0(x3_y16),
    .I1(x3_y17),
    .I2(x2_y20),
    .I3(x3_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010001100010)
) lut_6_20 (
    .O(x6_y20),
    .I0(1'b0),
    .I1(x3_y23),
    .I2(x3_y18),
    .I3(x3_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111001101100)
) lut_7_20 (
    .O(x7_y20),
    .I0(x5_y20),
    .I1(x5_y20),
    .I2(1'b0),
    .I3(x4_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110101000000)
) lut_8_20 (
    .O(x8_y20),
    .I0(x5_y15),
    .I1(1'b0),
    .I2(x6_y22),
    .I3(x5_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000011000000)
) lut_9_20 (
    .O(x9_y20),
    .I0(x7_y23),
    .I1(1'b0),
    .I2(x6_y22),
    .I3(x5_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011010100110)
) lut_10_20 (
    .O(x10_y20),
    .I0(x8_y16),
    .I1(x8_y19),
    .I2(x7_y20),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010000001011)
) lut_11_20 (
    .O(x11_y20),
    .I0(x9_y20),
    .I1(x8_y22),
    .I2(1'b0),
    .I3(x9_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001100100100)
) lut_12_20 (
    .O(x12_y20),
    .I0(x10_y17),
    .I1(x10_y19),
    .I2(x10_y20),
    .I3(x9_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001000010011)
) lut_13_20 (
    .O(x13_y20),
    .I0(x11_y23),
    .I1(1'b0),
    .I2(x11_y20),
    .I3(x11_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100110100011)
) lut_14_20 (
    .O(x14_y20),
    .I0(x12_y16),
    .I1(x12_y16),
    .I2(x12_y15),
    .I3(x11_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111000011010)
) lut_15_20 (
    .O(x15_y20),
    .I0(1'b0),
    .I1(x12_y24),
    .I2(x13_y21),
    .I3(x12_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111100100011)
) lut_16_20 (
    .O(x16_y20),
    .I0(x13_y19),
    .I1(x14_y20),
    .I2(x13_y24),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001111001110)
) lut_17_20 (
    .O(x17_y20),
    .I0(x14_y23),
    .I1(1'b0),
    .I2(x14_y24),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100000001011)
) lut_18_20 (
    .O(x18_y20),
    .I0(1'b0),
    .I1(x15_y25),
    .I2(x16_y21),
    .I3(x16_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011101010100)
) lut_19_20 (
    .O(x19_y20),
    .I0(x17_y17),
    .I1(x17_y17),
    .I2(x17_y22),
    .I3(x16_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101000101011)
) lut_20_20 (
    .O(x20_y20),
    .I0(1'b0),
    .I1(x18_y24),
    .I2(1'b0),
    .I3(x18_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000110001001)
) lut_21_20 (
    .O(x21_y20),
    .I0(1'b0),
    .I1(x18_y16),
    .I2(1'b0),
    .I3(x18_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111111100011)
) lut_22_20 (
    .O(x22_y20),
    .I0(1'b0),
    .I1(x19_y17),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101100010101)
) lut_23_20 (
    .O(x23_y20),
    .I0(x20_y16),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x21_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101011000100)
) lut_24_20 (
    .O(x24_y20),
    .I0(x22_y17),
    .I1(x21_y23),
    .I2(x22_y17),
    .I3(x22_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100000011001)
) lut_25_20 (
    .O(x25_y20),
    .I0(x23_y23),
    .I1(x23_y18),
    .I2(x23_y22),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110001001000)
) lut_26_20 (
    .O(x26_y20),
    .I0(x24_y16),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x24_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111011100001)
) lut_27_20 (
    .O(x27_y20),
    .I0(x25_y20),
    .I1(x25_y18),
    .I2(x25_y21),
    .I3(x24_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000101101110)
) lut_28_20 (
    .O(x28_y20),
    .I0(x25_y21),
    .I1(x25_y24),
    .I2(x26_y20),
    .I3(x26_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001010100110)
) lut_29_20 (
    .O(x29_y20),
    .I0(x27_y25),
    .I1(x27_y24),
    .I2(x27_y17),
    .I3(x26_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001010110101)
) lut_30_20 (
    .O(x30_y20),
    .I0(x28_y18),
    .I1(x27_y15),
    .I2(x28_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101100001000)
) lut_31_20 (
    .O(x31_y20),
    .I0(1'b0),
    .I1(x28_y20),
    .I2(x29_y18),
    .I3(x28_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010010111010)
) lut_32_20 (
    .O(x32_y20),
    .I0(x30_y22),
    .I1(x29_y17),
    .I2(x30_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100011001100)
) lut_33_20 (
    .O(x33_y20),
    .I0(x31_y16),
    .I1(x30_y23),
    .I2(x30_y15),
    .I3(x30_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011000001000)
) lut_34_20 (
    .O(x34_y20),
    .I0(x32_y17),
    .I1(x31_y16),
    .I2(1'b0),
    .I3(x32_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011001111110)
) lut_35_20 (
    .O(x35_y20),
    .I0(x32_y25),
    .I1(x32_y20),
    .I2(x32_y18),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110000010010)
) lut_36_20 (
    .O(x36_y20),
    .I0(x34_y21),
    .I1(x34_y15),
    .I2(x34_y17),
    .I3(x33_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101100000001)
) lut_37_20 (
    .O(x37_y20),
    .I0(1'b0),
    .I1(x34_y20),
    .I2(x34_y21),
    .I3(x34_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010010110000)
) lut_38_20 (
    .O(x38_y20),
    .I0(x36_y20),
    .I1(x35_y25),
    .I2(x35_y15),
    .I3(x35_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100010001111)
) lut_39_20 (
    .O(x39_y20),
    .I0(x37_y24),
    .I1(x37_y24),
    .I2(x36_y23),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110001110101)
) lut_40_20 (
    .O(x40_y20),
    .I0(x37_y24),
    .I1(x38_y15),
    .I2(x37_y20),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101100010110)
) lut_41_20 (
    .O(x41_y20),
    .I0(x39_y17),
    .I1(x38_y22),
    .I2(1'b0),
    .I3(x39_y15)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110001111100)
) lut_42_20 (
    .O(x42_y20),
    .I0(1'b0),
    .I1(x40_y25),
    .I2(x39_y25),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011001010000)
) lut_43_20 (
    .O(x43_y20),
    .I0(x40_y25),
    .I1(x40_y25),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101000111000)
) lut_44_20 (
    .O(x44_y20),
    .I0(x42_y17),
    .I1(x42_y21),
    .I2(1'b0),
    .I3(x41_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010001101011)
) lut_45_20 (
    .O(x45_y20),
    .I0(x42_y23),
    .I1(1'b0),
    .I2(x43_y17),
    .I3(x43_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001100000011)
) lut_46_20 (
    .O(x46_y20),
    .I0(1'b0),
    .I1(x43_y18),
    .I2(1'b0),
    .I3(x43_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101100101111)
) lut_47_20 (
    .O(x47_y20),
    .I0(x44_y21),
    .I1(x44_y25),
    .I2(x45_y23),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100011101101)
) lut_48_20 (
    .O(x48_y20),
    .I0(1'b0),
    .I1(x45_y20),
    .I2(x46_y19),
    .I3(x46_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100011000111)
) lut_49_20 (
    .O(x49_y20),
    .I0(x47_y22),
    .I1(x47_y24),
    .I2(x47_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011110010011)
) lut_50_20 (
    .O(x50_y20),
    .I0(x48_y20),
    .I1(x47_y16),
    .I2(x48_y23),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001111111101)
) lut_51_20 (
    .O(x51_y20),
    .I0(x48_y16),
    .I1(x49_y16),
    .I2(x48_y23),
    .I3(x49_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000000101001)
) lut_52_20 (
    .O(x52_y20),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x49_y16),
    .I3(x49_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110001000111)
) lut_53_20 (
    .O(x53_y20),
    .I0(x51_y24),
    .I1(x50_y20),
    .I2(1'b0),
    .I3(x51_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011110101111)
) lut_54_20 (
    .O(x54_y20),
    .I0(1'b0),
    .I1(x52_y17),
    .I2(x52_y24),
    .I3(x51_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111110101011)
) lut_55_20 (
    .O(x55_y20),
    .I0(x53_y23),
    .I1(x52_y15),
    .I2(x53_y20),
    .I3(x53_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000011101111)
) lut_56_20 (
    .O(x56_y20),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x53_y17),
    .I3(x53_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011000000011)
) lut_57_20 (
    .O(x57_y20),
    .I0(x54_y15),
    .I1(x54_y22),
    .I2(1'b0),
    .I3(x54_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010000100001)
) lut_58_20 (
    .O(x58_y20),
    .I0(1'b0),
    .I1(x56_y20),
    .I2(x55_y23),
    .I3(x56_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101010110011)
) lut_59_20 (
    .O(x59_y20),
    .I0(x56_y17),
    .I1(x56_y24),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111101010001)
) lut_60_20 (
    .O(x60_y20),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x58_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100010110111)
) lut_61_20 (
    .O(x61_y20),
    .I0(x58_y18),
    .I1(x58_y22),
    .I2(1'b0),
    .I3(x59_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011010000011)
) lut_62_20 (
    .O(x62_y20),
    .I0(x59_y16),
    .I1(1'b0),
    .I2(x60_y22),
    .I3(x59_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011001000111)
) lut_0_21 (
    .O(x0_y21),
    .I0(in2),
    .I1(in5),
    .I2(in8),
    .I3(in3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110100001000)
) lut_1_21 (
    .O(x1_y21),
    .I0(1'b0),
    .I1(in1),
    .I2(in2),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000001100100)
) lut_2_21 (
    .O(x2_y21),
    .I0(in2),
    .I1(1'b0),
    .I2(in1),
    .I3(in3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111101110100)
) lut_3_21 (
    .O(x3_y21),
    .I0(in1),
    .I1(x1_y26),
    .I2(1'b0),
    .I3(in5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000001000000)
) lut_4_21 (
    .O(x4_y21),
    .I0(x2_y17),
    .I1(x1_y22),
    .I2(1'b0),
    .I3(x1_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111100111101)
) lut_5_21 (
    .O(x5_y21),
    .I0(x2_y26),
    .I1(x3_y16),
    .I2(x3_y17),
    .I3(x3_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101101001010)
) lut_6_21 (
    .O(x6_y21),
    .I0(x4_y17),
    .I1(1'b0),
    .I2(x3_y17),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001101011101)
) lut_7_21 (
    .O(x7_y21),
    .I0(x4_y16),
    .I1(x5_y26),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001001001100)
) lut_8_21 (
    .O(x8_y21),
    .I0(x5_y20),
    .I1(x6_y24),
    .I2(x6_y20),
    .I3(x5_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100110101001)
) lut_9_21 (
    .O(x9_y21),
    .I0(x7_y19),
    .I1(x6_y18),
    .I2(x6_y20),
    .I3(x5_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101000011011)
) lut_10_21 (
    .O(x10_y21),
    .I0(1'b0),
    .I1(x8_y18),
    .I2(x7_y16),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010001101001)
) lut_11_21 (
    .O(x11_y21),
    .I0(1'b0),
    .I1(x9_y22),
    .I2(1'b0),
    .I3(x9_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111000110100)
) lut_12_21 (
    .O(x12_y21),
    .I0(x10_y22),
    .I1(x9_y21),
    .I2(1'b0),
    .I3(x9_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010011010010)
) lut_13_21 (
    .O(x13_y21),
    .I0(x10_y16),
    .I1(1'b0),
    .I2(x11_y17),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000000000000)
) lut_14_21 (
    .O(x14_y21),
    .I0(x11_y19),
    .I1(x12_y26),
    .I2(1'b0),
    .I3(x11_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111101000110)
) lut_15_21 (
    .O(x15_y21),
    .I0(x13_y21),
    .I1(1'b0),
    .I2(x13_y20),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110101101011)
) lut_16_21 (
    .O(x16_y21),
    .I0(x13_y20),
    .I1(x13_y20),
    .I2(x13_y24),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110000011110)
) lut_17_21 (
    .O(x17_y21),
    .I0(x15_y18),
    .I1(x15_y17),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001100001101)
) lut_18_21 (
    .O(x18_y21),
    .I0(x15_y24),
    .I1(x16_y19),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011100011010)
) lut_19_21 (
    .O(x19_y21),
    .I0(x16_y25),
    .I1(x16_y26),
    .I2(x17_y22),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101001010000)
) lut_20_21 (
    .O(x20_y21),
    .I0(x18_y25),
    .I1(1'b0),
    .I2(x18_y22),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000110010100)
) lut_21_21 (
    .O(x21_y21),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x18_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001111001100)
) lut_22_21 (
    .O(x22_y21),
    .I0(x20_y19),
    .I1(x20_y19),
    .I2(x20_y21),
    .I3(x19_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111011000010)
) lut_23_21 (
    .O(x23_y21),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x20_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100110111000)
) lut_24_21 (
    .O(x24_y21),
    .I0(1'b0),
    .I1(x21_y21),
    .I2(x21_y22),
    .I3(x21_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000100110100)
) lut_25_21 (
    .O(x25_y21),
    .I0(x23_y24),
    .I1(x22_y22),
    .I2(x23_y20),
    .I3(x22_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011110011110)
) lut_26_21 (
    .O(x26_y21),
    .I0(x23_y23),
    .I1(1'b0),
    .I2(x24_y19),
    .I3(x23_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010010000100)
) lut_27_21 (
    .O(x27_y21),
    .I0(x25_y24),
    .I1(1'b0),
    .I2(x25_y26),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001101001010)
) lut_28_21 (
    .O(x28_y21),
    .I0(x25_y24),
    .I1(x25_y17),
    .I2(1'b0),
    .I3(x26_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000011010111)
) lut_29_21 (
    .O(x29_y21),
    .I0(x27_y20),
    .I1(x27_y21),
    .I2(x27_y18),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000010010000)
) lut_30_21 (
    .O(x30_y21),
    .I0(x27_y18),
    .I1(x27_y24),
    .I2(x28_y21),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100001010101)
) lut_31_21 (
    .O(x31_y21),
    .I0(x29_y26),
    .I1(x29_y26),
    .I2(x29_y24),
    .I3(x29_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000110110111)
) lut_32_21 (
    .O(x32_y21),
    .I0(x30_y24),
    .I1(x29_y22),
    .I2(x29_y26),
    .I3(x30_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001010110001)
) lut_33_21 (
    .O(x33_y21),
    .I0(1'b0),
    .I1(x31_y16),
    .I2(x31_y25),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001100110100)
) lut_34_21 (
    .O(x34_y21),
    .I0(x32_y26),
    .I1(x31_y25),
    .I2(x31_y17),
    .I3(x32_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101001101001)
) lut_35_21 (
    .O(x35_y21),
    .I0(x32_y17),
    .I1(x32_y23),
    .I2(x32_y26),
    .I3(x32_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100100100110)
) lut_36_21 (
    .O(x36_y21),
    .I0(x33_y18),
    .I1(x34_y16),
    .I2(x34_y22),
    .I3(x33_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001100101101)
) lut_37_21 (
    .O(x37_y21),
    .I0(x34_y25),
    .I1(x34_y16),
    .I2(1'b0),
    .I3(x34_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101110110101)
) lut_38_21 (
    .O(x38_y21),
    .I0(x35_y19),
    .I1(x35_y19),
    .I2(x35_y20),
    .I3(x36_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100100101100)
) lut_39_21 (
    .O(x39_y21),
    .I0(x36_y19),
    .I1(x36_y20),
    .I2(1'b0),
    .I3(x37_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000101110101)
) lut_40_21 (
    .O(x40_y21),
    .I0(x37_y18),
    .I1(x38_y23),
    .I2(x37_y20),
    .I3(x37_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100111111001)
) lut_41_21 (
    .O(x41_y21),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x39_y20),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010111110101)
) lut_42_21 (
    .O(x42_y21),
    .I0(1'b0),
    .I1(x40_y22),
    .I2(x39_y21),
    .I3(x39_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011110010100)
) lut_43_21 (
    .O(x43_y21),
    .I0(x40_y24),
    .I1(1'b0),
    .I2(x41_y20),
    .I3(x41_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000100110001)
) lut_44_21 (
    .O(x44_y21),
    .I0(x41_y17),
    .I1(1'b0),
    .I2(x42_y22),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111100111100)
) lut_45_21 (
    .O(x45_y21),
    .I0(x42_y17),
    .I1(x42_y26),
    .I2(x43_y23),
    .I3(x42_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101100111000)
) lut_46_21 (
    .O(x46_y21),
    .I0(x44_y22),
    .I1(x44_y18),
    .I2(x43_y22),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011110010010)
) lut_47_21 (
    .O(x47_y21),
    .I0(1'b0),
    .I1(x44_y22),
    .I2(x44_y19),
    .I3(x44_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111000110010)
) lut_48_21 (
    .O(x48_y21),
    .I0(1'b0),
    .I1(x45_y23),
    .I2(1'b0),
    .I3(x45_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111100110101)
) lut_49_21 (
    .O(x49_y21),
    .I0(x47_y24),
    .I1(x46_y19),
    .I2(x47_y21),
    .I3(x46_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110001111110)
) lut_50_21 (
    .O(x50_y21),
    .I0(x48_y19),
    .I1(1'b0),
    .I2(x47_y19),
    .I3(x48_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100111001010)
) lut_51_21 (
    .O(x51_y21),
    .I0(1'b0),
    .I1(x48_y16),
    .I2(x49_y16),
    .I3(x49_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010010011000)
) lut_52_21 (
    .O(x52_y21),
    .I0(x50_y18),
    .I1(x49_y16),
    .I2(x49_y18),
    .I3(x50_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111011000110)
) lut_53_21 (
    .O(x53_y21),
    .I0(x50_y16),
    .I1(x51_y16),
    .I2(x51_y18),
    .I3(x51_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101110110010)
) lut_54_21 (
    .O(x54_y21),
    .I0(x51_y21),
    .I1(x52_y22),
    .I2(1'b0),
    .I3(x52_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100010110101)
) lut_55_21 (
    .O(x55_y21),
    .I0(1'b0),
    .I1(x53_y22),
    .I2(x53_y23),
    .I3(x53_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000111111100)
) lut_56_21 (
    .O(x56_y21),
    .I0(x53_y19),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x53_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101100110001)
) lut_57_21 (
    .O(x57_y21),
    .I0(x54_y22),
    .I1(1'b0),
    .I2(x55_y25),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101000111001)
) lut_58_21 (
    .O(x58_y21),
    .I0(x55_y21),
    .I1(x56_y22),
    .I2(x55_y22),
    .I3(x55_y16)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111010100010)
) lut_59_21 (
    .O(x59_y21),
    .I0(x57_y20),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x56_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111010111110)
) lut_60_21 (
    .O(x60_y21),
    .I0(x58_y17),
    .I1(x57_y20),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011111011001)
) lut_61_21 (
    .O(x61_y21),
    .I0(x59_y23),
    .I1(x59_y17),
    .I2(x58_y25),
    .I3(x59_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111001010011)
) lut_62_21 (
    .O(x62_y21),
    .I0(x59_y17),
    .I1(1'b0),
    .I2(x60_y26),
    .I3(x59_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110101010010)
) lut_0_22 (
    .O(x0_y22),
    .I0(1'b0),
    .I1(in5),
    .I2(1'b0),
    .I3(in3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100110010110)
) lut_1_22 (
    .O(x1_y22),
    .I0(1'b0),
    .I1(in9),
    .I2(in7),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000001010110)
) lut_2_22 (
    .O(x2_y22),
    .I0(in3),
    .I1(1'b0),
    .I2(in5),
    .I3(in5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000101100011)
) lut_3_22 (
    .O(x3_y22),
    .I0(in4),
    .I1(1'b0),
    .I2(in8),
    .I3(x1_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001001011100)
) lut_4_22 (
    .O(x4_y22),
    .I0(1'b0),
    .I1(x1_y19),
    .I2(x1_y21),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100111100000)
) lut_5_22 (
    .O(x5_y22),
    .I0(x3_y20),
    .I1(1'b0),
    .I2(x2_y23),
    .I3(x2_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000100011101)
) lut_6_22 (
    .O(x6_y22),
    .I0(x3_y24),
    .I1(x3_y23),
    .I2(x3_y24),
    .I3(x4_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000011000010)
) lut_7_22 (
    .O(x7_y22),
    .I0(x4_y17),
    .I1(x5_y18),
    .I2(x4_y21),
    .I3(x4_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001110111110)
) lut_8_22 (
    .O(x8_y22),
    .I0(x5_y18),
    .I1(x6_y24),
    .I2(1'b0),
    .I3(x6_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011011100110)
) lut_9_22 (
    .O(x9_y22),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x6_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010000011111)
) lut_10_22 (
    .O(x10_y22),
    .I0(x7_y22),
    .I1(x7_y19),
    .I2(x8_y17),
    .I3(x8_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101101000100)
) lut_11_22 (
    .O(x11_y22),
    .I0(x9_y17),
    .I1(x8_y26),
    .I2(x8_y23),
    .I3(x9_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000111011100)
) lut_12_22 (
    .O(x12_y22),
    .I0(1'b0),
    .I1(x10_y25),
    .I2(x9_y18),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110111000100)
) lut_13_22 (
    .O(x13_y22),
    .I0(x11_y24),
    .I1(x11_y25),
    .I2(x11_y18),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010010100110)
) lut_14_22 (
    .O(x14_y22),
    .I0(x12_y19),
    .I1(1'b0),
    .I2(x11_y17),
    .I3(x12_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101010011011)
) lut_15_22 (
    .O(x15_y22),
    .I0(x12_y25),
    .I1(1'b0),
    .I2(x12_y20),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010100110110)
) lut_16_22 (
    .O(x16_y22),
    .I0(1'b0),
    .I1(x14_y17),
    .I2(1'b0),
    .I3(x14_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101100101111)
) lut_17_22 (
    .O(x17_y22),
    .I0(x14_y20),
    .I1(x14_y21),
    .I2(x14_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011010001100)
) lut_18_22 (
    .O(x18_y22),
    .I0(x16_y23),
    .I1(x16_y27),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101111000010)
) lut_19_22 (
    .O(x19_y22),
    .I0(x16_y22),
    .I1(x16_y18),
    .I2(x16_y22),
    .I3(x16_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101101111011)
) lut_20_22 (
    .O(x20_y22),
    .I0(1'b0),
    .I1(x17_y18),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000101110000)
) lut_21_22 (
    .O(x21_y22),
    .I0(1'b0),
    .I1(x18_y22),
    .I2(1'b0),
    .I3(x18_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100001111100)
) lut_22_22 (
    .O(x22_y22),
    .I0(x19_y17),
    .I1(x20_y20),
    .I2(x19_y17),
    .I3(x19_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111111001010)
) lut_23_22 (
    .O(x23_y22),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x20_y25),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000001110001)
) lut_24_22 (
    .O(x24_y22),
    .I0(x21_y24),
    .I1(x21_y18),
    .I2(x22_y22),
    .I3(x21_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001111010011)
) lut_25_22 (
    .O(x25_y22),
    .I0(1'b0),
    .I1(x22_y24),
    .I2(x23_y18),
    .I3(x23_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011100001010)
) lut_26_22 (
    .O(x26_y22),
    .I0(1'b0),
    .I1(x23_y20),
    .I2(x23_y19),
    .I3(x23_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001010010100)
) lut_27_22 (
    .O(x27_y22),
    .I0(x24_y21),
    .I1(x25_y21),
    .I2(1'b0),
    .I3(x24_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011101100000)
) lut_28_22 (
    .O(x28_y22),
    .I0(x25_y21),
    .I1(x25_y26),
    .I2(x26_y24),
    .I3(x25_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111001110010)
) lut_29_22 (
    .O(x29_y22),
    .I0(x27_y21),
    .I1(x27_y19),
    .I2(x27_y17),
    .I3(x27_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001110101101)
) lut_30_22 (
    .O(x30_y22),
    .I0(1'b0),
    .I1(x28_y20),
    .I2(x27_y20),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100101111111)
) lut_31_22 (
    .O(x31_y22),
    .I0(1'b0),
    .I1(x29_y23),
    .I2(1'b0),
    .I3(x29_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000101010111)
) lut_32_22 (
    .O(x32_y22),
    .I0(x29_y26),
    .I1(x29_y27),
    .I2(x29_y26),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001000111011)
) lut_33_22 (
    .O(x33_y22),
    .I0(x31_y23),
    .I1(x31_y26),
    .I2(x31_y19),
    .I3(x31_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110000010001)
) lut_34_22 (
    .O(x34_y22),
    .I0(x32_y24),
    .I1(x31_y25),
    .I2(x31_y22),
    .I3(x32_y17)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110010101100)
) lut_35_22 (
    .O(x35_y22),
    .I0(x32_y24),
    .I1(x33_y27),
    .I2(x32_y24),
    .I3(x32_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000101101010)
) lut_36_22 (
    .O(x36_y22),
    .I0(x33_y23),
    .I1(x33_y21),
    .I2(x33_y23),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101001011001)
) lut_37_22 (
    .O(x37_y22),
    .I0(x35_y20),
    .I1(x34_y17),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001110000110)
) lut_38_22 (
    .O(x38_y22),
    .I0(x36_y27),
    .I1(x36_y21),
    .I2(x36_y21),
    .I3(x35_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001100000011)
) lut_39_22 (
    .O(x39_y22),
    .I0(1'b0),
    .I1(x37_y27),
    .I2(x36_y22),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011010100001)
) lut_40_22 (
    .O(x40_y22),
    .I0(x37_y27),
    .I1(x38_y19),
    .I2(x38_y21),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111100111010)
) lut_41_22 (
    .O(x41_y22),
    .I0(1'b0),
    .I1(x38_y26),
    .I2(x39_y26),
    .I3(x39_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000011000101)
) lut_42_22 (
    .O(x42_y22),
    .I0(1'b0),
    .I1(x39_y21),
    .I2(x40_y21),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001010010101)
) lut_43_22 (
    .O(x43_y22),
    .I0(x41_y21),
    .I1(x41_y18),
    .I2(1'b0),
    .I3(x40_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101001110100)
) lut_44_22 (
    .O(x44_y22),
    .I0(x42_y17),
    .I1(x42_y21),
    .I2(x41_y20),
    .I3(x41_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111101111010)
) lut_45_22 (
    .O(x45_y22),
    .I0(x42_y20),
    .I1(x43_y22),
    .I2(x43_y23),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000011001100)
) lut_46_22 (
    .O(x46_y22),
    .I0(x43_y26),
    .I1(1'b0),
    .I2(x44_y20),
    .I3(x43_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000001001011)
) lut_47_22 (
    .O(x47_y22),
    .I0(x44_y21),
    .I1(x45_y19),
    .I2(x45_y17),
    .I3(x45_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101010100000)
) lut_48_22 (
    .O(x48_y22),
    .I0(x46_y22),
    .I1(x46_y25),
    .I2(1'b0),
    .I3(x46_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001101101101)
) lut_49_22 (
    .O(x49_y22),
    .I0(1'b0),
    .I1(x46_y18),
    .I2(x47_y25),
    .I3(x46_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001010001011)
) lut_50_22 (
    .O(x50_y22),
    .I0(1'b0),
    .I1(x48_y17),
    .I2(1'b0),
    .I3(x48_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100010010100)
) lut_51_22 (
    .O(x51_y22),
    .I0(1'b0),
    .I1(x49_y18),
    .I2(x49_y25),
    .I3(x49_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111001111000)
) lut_52_22 (
    .O(x52_y22),
    .I0(x50_y19),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001000101000)
) lut_53_22 (
    .O(x53_y22),
    .I0(x50_y24),
    .I1(1'b0),
    .I2(x51_y25),
    .I3(x50_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000010100100)
) lut_54_22 (
    .O(x54_y22),
    .I0(x52_y25),
    .I1(x51_y26),
    .I2(x52_y19),
    .I3(x51_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101011100101)
) lut_55_22 (
    .O(x55_y22),
    .I0(x53_y27),
    .I1(x52_y18),
    .I2(x53_y26),
    .I3(x53_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000101110101)
) lut_56_22 (
    .O(x56_y22),
    .I0(x53_y20),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x53_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100110111000)
) lut_57_22 (
    .O(x57_y22),
    .I0(x55_y19),
    .I1(x55_y26),
    .I2(1'b0),
    .I3(x55_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110000110101)
) lut_58_22 (
    .O(x58_y22),
    .I0(x56_y18),
    .I1(x56_y23),
    .I2(x55_y20),
    .I3(x56_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001001011110)
) lut_59_22 (
    .O(x59_y22),
    .I0(x57_y27),
    .I1(x57_y19),
    .I2(1'b0),
    .I3(x57_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000110111000)
) lut_60_22 (
    .O(x60_y22),
    .I0(x58_y24),
    .I1(x57_y27),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011001110011)
) lut_61_22 (
    .O(x61_y22),
    .I0(x59_y20),
    .I1(x59_y17),
    .I2(1'b0),
    .I3(x59_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010101010010)
) lut_62_22 (
    .O(x62_y22),
    .I0(x60_y19),
    .I1(x60_y17),
    .I2(1'b0),
    .I3(x59_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011111101110)
) lut_0_23 (
    .O(x0_y23),
    .I0(1'b0),
    .I1(1'b0),
    .I2(in4),
    .I3(in3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101001101101)
) lut_1_23 (
    .O(x1_y23),
    .I0(in2),
    .I1(in1),
    .I2(in1),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110110000011)
) lut_2_23 (
    .O(x2_y23),
    .I0(1'b0),
    .I1(in3),
    .I2(1'b0),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010001001000)
) lut_3_23 (
    .O(x3_y23),
    .I0(x1_y20),
    .I1(x1_y25),
    .I2(in0),
    .I3(x1_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001100100000)
) lut_4_23 (
    .O(x4_y23),
    .I0(x1_y27),
    .I1(x2_y27),
    .I2(x2_y21),
    .I3(x2_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111101101100)
) lut_5_23 (
    .O(x5_y23),
    .I0(1'b0),
    .I1(x3_y24),
    .I2(x2_y21),
    .I3(x2_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101100000110)
) lut_6_23 (
    .O(x6_y23),
    .I0(x3_y22),
    .I1(1'b0),
    .I2(x4_y28),
    .I3(x3_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011110001000)
) lut_7_23 (
    .O(x7_y23),
    .I0(x4_y19),
    .I1(1'b0),
    .I2(x4_y22),
    .I3(x4_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011001100010)
) lut_8_23 (
    .O(x8_y23),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x5_y23),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000101100000)
) lut_9_23 (
    .O(x9_y23),
    .I0(x7_y22),
    .I1(1'b0),
    .I2(x5_y23),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010111100100)
) lut_10_23 (
    .O(x10_y23),
    .I0(x8_y21),
    .I1(x8_y27),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110000111001)
) lut_11_23 (
    .O(x11_y23),
    .I0(x9_y20),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x8_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011110111101)
) lut_12_23 (
    .O(x12_y23),
    .I0(x10_y28),
    .I1(x9_y19),
    .I2(1'b0),
    .I3(x10_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011101010011)
) lut_13_23 (
    .O(x13_y23),
    .I0(x10_y25),
    .I1(x11_y19),
    .I2(1'b0),
    .I3(x10_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100110001001)
) lut_14_23 (
    .O(x14_y23),
    .I0(x12_y25),
    .I1(x11_y27),
    .I2(x12_y23),
    .I3(x11_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001101100011)
) lut_15_23 (
    .O(x15_y23),
    .I0(x13_y28),
    .I1(x13_y23),
    .I2(x13_y21),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000001001100)
) lut_16_23 (
    .O(x16_y23),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x13_y20),
    .I3(x13_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011101101001)
) lut_17_23 (
    .O(x17_y23),
    .I0(x15_y21),
    .I1(x14_y24),
    .I2(1'b0),
    .I3(x14_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010100011100)
) lut_18_23 (
    .O(x18_y23),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x16_y20),
    .I3(x15_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001011100100)
) lut_19_23 (
    .O(x19_y23),
    .I0(x16_y25),
    .I1(x17_y23),
    .I2(x16_y22),
    .I3(x17_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101111101001)
) lut_20_23 (
    .O(x20_y23),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110110000110)
) lut_21_23 (
    .O(x21_y23),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x19_y25),
    .I3(x18_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100110100111)
) lut_22_23 (
    .O(x22_y23),
    .I0(x19_y26),
    .I1(x20_y27),
    .I2(x19_y20),
    .I3(x20_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001000101111)
) lut_23_23 (
    .O(x23_y23),
    .I0(x21_y18),
    .I1(1'b0),
    .I2(x21_y26),
    .I3(x20_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000011011110)
) lut_24_23 (
    .O(x24_y23),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x21_y25),
    .I3(x22_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111000111011)
) lut_25_23 (
    .O(x25_y23),
    .I0(x22_y26),
    .I1(x22_y19),
    .I2(x22_y23),
    .I3(x22_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100010101110)
) lut_26_23 (
    .O(x26_y23),
    .I0(x24_y25),
    .I1(x24_y21),
    .I2(x24_y19),
    .I3(x24_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111101011110)
) lut_27_23 (
    .O(x27_y23),
    .I0(x24_y27),
    .I1(x24_y19),
    .I2(x25_y24),
    .I3(x24_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101101110111)
) lut_28_23 (
    .O(x28_y23),
    .I0(x26_y27),
    .I1(1'b0),
    .I2(x25_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101100110011)
) lut_29_23 (
    .O(x29_y23),
    .I0(x26_y19),
    .I1(x26_y24),
    .I2(x27_y26),
    .I3(x26_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000110101001)
) lut_30_23 (
    .O(x30_y23),
    .I0(1'b0),
    .I1(x27_y27),
    .I2(1'b0),
    .I3(x27_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110010100001)
) lut_31_23 (
    .O(x31_y23),
    .I0(x29_y20),
    .I1(1'b0),
    .I2(x29_y28),
    .I3(x28_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011001101100)
) lut_32_23 (
    .O(x32_y23),
    .I0(x29_y19),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x29_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101010000011)
) lut_33_23 (
    .O(x33_y23),
    .I0(x30_y27),
    .I1(x31_y18),
    .I2(x31_y22),
    .I3(x31_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111001110101)
) lut_34_23 (
    .O(x34_y23),
    .I0(x32_y28),
    .I1(1'b0),
    .I2(x31_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101011110111)
) lut_35_23 (
    .O(x35_y23),
    .I0(x33_y19),
    .I1(x32_y20),
    .I2(1'b0),
    .I3(x32_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100110001011)
) lut_36_23 (
    .O(x36_y23),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x33_y23),
    .I3(x34_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110001110110)
) lut_37_23 (
    .O(x37_y23),
    .I0(x34_y26),
    .I1(x34_y21),
    .I2(x34_y27),
    .I3(x34_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101110100111)
) lut_38_23 (
    .O(x38_y23),
    .I0(1'b0),
    .I1(x35_y25),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011101000000)
) lut_39_23 (
    .O(x39_y23),
    .I0(1'b0),
    .I1(x37_y20),
    .I2(x37_y19),
    .I3(x36_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010111000100)
) lut_40_23 (
    .O(x40_y23),
    .I0(1'b0),
    .I1(x38_y26),
    .I2(x37_y25),
    .I3(x38_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111100111000)
) lut_41_23 (
    .O(x41_y23),
    .I0(x38_y19),
    .I1(x39_y24),
    .I2(x39_y20),
    .I3(x39_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111010100010)
) lut_42_23 (
    .O(x42_y23),
    .I0(x39_y26),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x39_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001001011111)
) lut_43_23 (
    .O(x43_y23),
    .I0(x40_y19),
    .I1(x40_y25),
    .I2(x41_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010010010011)
) lut_44_23 (
    .O(x44_y23),
    .I0(1'b0),
    .I1(x42_y26),
    .I2(x42_y20),
    .I3(x41_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100111000100)
) lut_45_23 (
    .O(x45_y23),
    .I0(1'b0),
    .I1(x42_y27),
    .I2(x43_y25),
    .I3(x42_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101111010010)
) lut_46_23 (
    .O(x46_y23),
    .I0(x43_y19),
    .I1(x44_y24),
    .I2(x44_y21),
    .I3(x43_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011000101001)
) lut_47_23 (
    .O(x47_y23),
    .I0(x44_y19),
    .I1(1'b0),
    .I2(x44_y21),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000010011010)
) lut_48_23 (
    .O(x48_y23),
    .I0(x45_y19),
    .I1(x46_y22),
    .I2(1'b0),
    .I3(x45_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000101000111)
) lut_49_23 (
    .O(x49_y23),
    .I0(x47_y25),
    .I1(x47_y21),
    .I2(x46_y23),
    .I3(x46_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100111000110)
) lut_50_23 (
    .O(x50_y23),
    .I0(x48_y27),
    .I1(x48_y22),
    .I2(x48_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000011101100)
) lut_51_23 (
    .O(x51_y23),
    .I0(x48_y19),
    .I1(x48_y25),
    .I2(x48_y19),
    .I3(x49_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000001000100)
) lut_52_23 (
    .O(x52_y23),
    .I0(x50_y18),
    .I1(x50_y23),
    .I2(1'b0),
    .I3(x50_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010110010100)
) lut_53_23 (
    .O(x53_y23),
    .I0(1'b0),
    .I1(x50_y18),
    .I2(1'b0),
    .I3(x50_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100100001010)
) lut_54_23 (
    .O(x54_y23),
    .I0(x51_y24),
    .I1(x52_y22),
    .I2(x51_y28),
    .I3(x51_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011000111100)
) lut_55_23 (
    .O(x55_y23),
    .I0(x53_y20),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010011100000)
) lut_56_23 (
    .O(x56_y23),
    .I0(x54_y24),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101000111110)
) lut_57_23 (
    .O(x57_y23),
    .I0(x54_y24),
    .I1(x54_y24),
    .I2(1'b0),
    .I3(x55_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010101001100)
) lut_58_23 (
    .O(x58_y23),
    .I0(x56_y18),
    .I1(1'b0),
    .I2(x55_y18),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011101001001)
) lut_59_23 (
    .O(x59_y23),
    .I0(x57_y22),
    .I1(x57_y23),
    .I2(x57_y25),
    .I3(x57_y18)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001001011001)
) lut_60_23 (
    .O(x60_y23),
    .I0(x58_y27),
    .I1(1'b0),
    .I2(x57_y20),
    .I3(x57_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100001001011)
) lut_61_23 (
    .O(x61_y23),
    .I0(x59_y22),
    .I1(x58_y22),
    .I2(x59_y18),
    .I3(x59_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101100110001)
) lut_62_23 (
    .O(x62_y23),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x59_y23),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100000110001)
) lut_0_24 (
    .O(x0_y24),
    .I0(1'b0),
    .I1(in1),
    .I2(1'b0),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110110000110)
) lut_1_24 (
    .O(x1_y24),
    .I0(in4),
    .I1(1'b0),
    .I2(in4),
    .I3(in5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001001011111)
) lut_2_24 (
    .O(x2_y24),
    .I0(in7),
    .I1(1'b0),
    .I2(in1),
    .I3(in1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011111111011)
) lut_3_24 (
    .O(x3_y24),
    .I0(1'b0),
    .I1(x1_y26),
    .I2(1'b0),
    .I3(x1_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000010001001)
) lut_4_24 (
    .O(x4_y24),
    .I0(x2_y25),
    .I1(x1_y22),
    .I2(x2_y24),
    .I3(x2_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000011000111)
) lut_5_24 (
    .O(x5_y24),
    .I0(x3_y19),
    .I1(1'b0),
    .I2(x3_y20),
    .I3(x2_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011000111110)
) lut_6_24 (
    .O(x6_y24),
    .I0(1'b0),
    .I1(x3_y23),
    .I2(1'b0),
    .I3(x4_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000101110011)
) lut_7_24 (
    .O(x7_y24),
    .I0(x5_y19),
    .I1(1'b0),
    .I2(x4_y22),
    .I3(x5_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110000100011)
) lut_8_24 (
    .O(x8_y24),
    .I0(x5_y22),
    .I1(x5_y24),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001000000010)
) lut_9_24 (
    .O(x9_y24),
    .I0(x6_y23),
    .I1(x6_y22),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110000101000)
) lut_10_24 (
    .O(x10_y24),
    .I0(x7_y23),
    .I1(x8_y26),
    .I2(x8_y20),
    .I3(x8_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000010010101)
) lut_11_24 (
    .O(x11_y24),
    .I0(x8_y21),
    .I1(1'b0),
    .I2(x9_y22),
    .I3(x9_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110011111010)
) lut_12_24 (
    .O(x12_y24),
    .I0(x10_y22),
    .I1(x10_y21),
    .I2(1'b0),
    .I3(x9_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010110000100)
) lut_13_24 (
    .O(x13_y24),
    .I0(x11_y22),
    .I1(x10_y26),
    .I2(x10_y25),
    .I3(x10_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010011001101)
) lut_14_24 (
    .O(x14_y24),
    .I0(x12_y26),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x11_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111011110000)
) lut_15_24 (
    .O(x15_y24),
    .I0(x13_y20),
    .I1(x13_y27),
    .I2(x13_y26),
    .I3(x12_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010111001010)
) lut_16_24 (
    .O(x16_y24),
    .I0(x14_y26),
    .I1(x13_y28),
    .I2(x14_y29),
    .I3(x14_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001001001010)
) lut_17_24 (
    .O(x17_y24),
    .I0(x14_y28),
    .I1(1'b0),
    .I2(x14_y21),
    .I3(x15_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101101010100)
) lut_18_24 (
    .O(x18_y24),
    .I0(x16_y23),
    .I1(x15_y29),
    .I2(x16_y25),
    .I3(x16_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011110000100)
) lut_19_24 (
    .O(x19_y24),
    .I0(x16_y24),
    .I1(x17_y22),
    .I2(x16_y28),
    .I3(x16_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101110001011)
) lut_20_24 (
    .O(x20_y24),
    .I0(x17_y27),
    .I1(x17_y27),
    .I2(x17_y27),
    .I3(x17_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010101010011)
) lut_21_24 (
    .O(x21_y24),
    .I0(x18_y24),
    .I1(1'b0),
    .I2(x19_y20),
    .I3(x18_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100011100000)
) lut_22_24 (
    .O(x22_y24),
    .I0(1'b0),
    .I1(x20_y22),
    .I2(x19_y29),
    .I3(x20_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010001111000)
) lut_23_24 (
    .O(x23_y24),
    .I0(x20_y22),
    .I1(x20_y22),
    .I2(x21_y20),
    .I3(x21_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101000100111)
) lut_24_24 (
    .O(x24_y24),
    .I0(x22_y24),
    .I1(x22_y20),
    .I2(x21_y25),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110101011000)
) lut_25_24 (
    .O(x25_y24),
    .I0(x23_y23),
    .I1(1'b0),
    .I2(x22_y25),
    .I3(x22_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101001111001)
) lut_26_24 (
    .O(x26_y24),
    .I0(x24_y21),
    .I1(1'b0),
    .I2(x23_y29),
    .I3(x23_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000011111001)
) lut_27_24 (
    .O(x27_y24),
    .I0(1'b0),
    .I1(x25_y20),
    .I2(x24_y26),
    .I3(x25_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011101000100)
) lut_28_24 (
    .O(x28_y24),
    .I0(x25_y20),
    .I1(1'b0),
    .I2(x25_y23),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011000011001)
) lut_29_24 (
    .O(x29_y24),
    .I0(x27_y19),
    .I1(x27_y21),
    .I2(1'b0),
    .I3(x27_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001011001011)
) lut_30_24 (
    .O(x30_y24),
    .I0(x28_y29),
    .I1(x28_y28),
    .I2(x28_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101101101101)
) lut_31_24 (
    .O(x31_y24),
    .I0(1'b0),
    .I1(x29_y19),
    .I2(x28_y22),
    .I3(x29_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001001011000)
) lut_32_24 (
    .O(x32_y24),
    .I0(1'b0),
    .I1(x30_y28),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000101100111)
) lut_33_24 (
    .O(x33_y24),
    .I0(x31_y19),
    .I1(1'b0),
    .I2(x31_y21),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110001111111)
) lut_34_24 (
    .O(x34_y24),
    .I0(1'b0),
    .I1(x31_y24),
    .I2(x31_y25),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100000011001)
) lut_35_24 (
    .O(x35_y24),
    .I0(x33_y20),
    .I1(x33_y19),
    .I2(x32_y21),
    .I3(x32_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100101111111)
) lut_36_24 (
    .O(x36_y24),
    .I0(x33_y29),
    .I1(x33_y29),
    .I2(x34_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111101101001)
) lut_37_24 (
    .O(x37_y24),
    .I0(x34_y29),
    .I1(x35_y27),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100010100011)
) lut_38_24 (
    .O(x38_y24),
    .I0(1'b0),
    .I1(x35_y25),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100101100100)
) lut_39_24 (
    .O(x39_y24),
    .I0(x37_y24),
    .I1(1'b0),
    .I2(x36_y27),
    .I3(x36_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111100000111)
) lut_40_24 (
    .O(x40_y24),
    .I0(x37_y26),
    .I1(1'b0),
    .I2(x37_y22),
    .I3(x38_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010011011010)
) lut_41_24 (
    .O(x41_y24),
    .I0(x39_y24),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x38_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010111010010)
) lut_42_24 (
    .O(x42_y24),
    .I0(x39_y22),
    .I1(x39_y27),
    .I2(x39_y24),
    .I3(x40_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000001010000)
) lut_43_24 (
    .O(x43_y24),
    .I0(x40_y20),
    .I1(1'b0),
    .I2(x41_y24),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111101001010)
) lut_44_24 (
    .O(x44_y24),
    .I0(x42_y22),
    .I1(x41_y21),
    .I2(x41_y22),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101101001011)
) lut_45_24 (
    .O(x45_y24),
    .I0(x42_y25),
    .I1(x43_y19),
    .I2(x43_y21),
    .I3(x43_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000110110101)
) lut_46_24 (
    .O(x46_y24),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x43_y21),
    .I3(x44_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101110001110)
) lut_47_24 (
    .O(x47_y24),
    .I0(x45_y26),
    .I1(x45_y19),
    .I2(x45_y24),
    .I3(x44_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100001101101)
) lut_48_24 (
    .O(x48_y24),
    .I0(1'b0),
    .I1(x46_y26),
    .I2(x45_y20),
    .I3(x46_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101001100101)
) lut_49_24 (
    .O(x49_y24),
    .I0(1'b0),
    .I1(x46_y20),
    .I2(x47_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111101010001)
) lut_50_24 (
    .O(x50_y24),
    .I0(x48_y26),
    .I1(x48_y26),
    .I2(x48_y21),
    .I3(x47_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101110011000)
) lut_51_24 (
    .O(x51_y24),
    .I0(x48_y19),
    .I1(x49_y25),
    .I2(x49_y29),
    .I3(x49_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000100011011)
) lut_52_24 (
    .O(x52_y24),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x50_y19)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000001101111)
) lut_53_24 (
    .O(x53_y24),
    .I0(1'b0),
    .I1(x50_y29),
    .I2(x51_y28),
    .I3(x51_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000100111100)
) lut_54_24 (
    .O(x54_y24),
    .I0(x52_y23),
    .I1(x52_y29),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010101110000)
) lut_55_24 (
    .O(x55_y24),
    .I0(1'b0),
    .I1(x52_y23),
    .I2(1'b0),
    .I3(x53_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100111000111)
) lut_56_24 (
    .O(x56_y24),
    .I0(x53_y23),
    .I1(x53_y19),
    .I2(1'b0),
    .I3(x53_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000100100100)
) lut_57_24 (
    .O(x57_y24),
    .I0(x55_y22),
    .I1(x55_y19),
    .I2(x54_y22),
    .I3(x54_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110110010110)
) lut_58_24 (
    .O(x58_y24),
    .I0(x56_y23),
    .I1(x56_y24),
    .I2(x55_y24),
    .I3(x55_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000000101001)
) lut_59_24 (
    .O(x59_y24),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x57_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010000000101)
) lut_60_24 (
    .O(x60_y24),
    .I0(x57_y28),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x58_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110100010101)
) lut_61_24 (
    .O(x61_y24),
    .I0(x58_y26),
    .I1(x59_y22),
    .I2(x59_y23),
    .I3(x59_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001011101110)
) lut_62_24 (
    .O(x62_y24),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x60_y20),
    .I3(x60_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101010011001)
) lut_0_25 (
    .O(x0_y25),
    .I0(in9),
    .I1(in6),
    .I2(in8),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110011000010)
) lut_1_25 (
    .O(x1_y25),
    .I0(in4),
    .I1(in1),
    .I2(in0),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001000100001)
) lut_2_25 (
    .O(x2_y25),
    .I0(in2),
    .I1(in0),
    .I2(1'b0),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100010010110)
) lut_3_25 (
    .O(x3_y25),
    .I0(in0),
    .I1(in6),
    .I2(in5),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110001011100)
) lut_4_25 (
    .O(x4_y25),
    .I0(1'b0),
    .I1(x1_y21),
    .I2(x1_y24),
    .I3(x2_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000100100100)
) lut_5_25 (
    .O(x5_y25),
    .I0(x3_y23),
    .I1(x3_y25),
    .I2(x2_y21),
    .I3(x2_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001111000011)
) lut_6_25 (
    .O(x6_y25),
    .I0(x4_y23),
    .I1(1'b0),
    .I2(x4_y25),
    .I3(x3_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000100111111)
) lut_7_25 (
    .O(x7_y25),
    .I0(x4_y23),
    .I1(x5_y22),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100011011001)
) lut_8_25 (
    .O(x8_y25),
    .I0(1'b0),
    .I1(x5_y23),
    .I2(x6_y27),
    .I3(x6_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011100001001)
) lut_9_25 (
    .O(x9_y25),
    .I0(x7_y30),
    .I1(x6_y24),
    .I2(x6_y27),
    .I3(x6_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001001001111)
) lut_10_25 (
    .O(x10_y25),
    .I0(1'b0),
    .I1(x8_y20),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001101111100)
) lut_11_25 (
    .O(x11_y25),
    .I0(x8_y25),
    .I1(x8_y29),
    .I2(x8_y23),
    .I3(x8_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001101001010)
) lut_12_25 (
    .O(x12_y25),
    .I0(1'b0),
    .I1(x10_y27),
    .I2(x9_y23),
    .I3(x10_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000001000010)
) lut_13_25 (
    .O(x13_y25),
    .I0(x10_y25),
    .I1(x10_y21),
    .I2(x10_y21),
    .I3(x11_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011111011010)
) lut_14_25 (
    .O(x14_y25),
    .I0(x11_y23),
    .I1(x12_y25),
    .I2(x12_y22),
    .I3(x12_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001100100111)
) lut_15_25 (
    .O(x15_y25),
    .I0(x13_y23),
    .I1(1'b0),
    .I2(x12_y21),
    .I3(x12_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000000010110)
) lut_16_25 (
    .O(x16_y25),
    .I0(1'b0),
    .I1(x14_y28),
    .I2(1'b0),
    .I3(x13_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111101011011)
) lut_17_25 (
    .O(x17_y25),
    .I0(x15_y25),
    .I1(x15_y22),
    .I2(x15_y22),
    .I3(x15_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110111110001)
) lut_18_25 (
    .O(x18_y25),
    .I0(1'b0),
    .I1(x15_y26),
    .I2(x15_y23),
    .I3(x15_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100010110011)
) lut_19_25 (
    .O(x19_y25),
    .I0(x16_y23),
    .I1(1'b0),
    .I2(x16_y23),
    .I3(x17_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100111010010)
) lut_20_25 (
    .O(x20_y25),
    .I0(x17_y28),
    .I1(1'b0),
    .I2(x18_y24),
    .I3(x17_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100100000111)
) lut_21_25 (
    .O(x21_y25),
    .I0(1'b0),
    .I1(x19_y30),
    .I2(1'b0),
    .I3(x18_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101110011000)
) lut_22_25 (
    .O(x22_y25),
    .I0(x19_y20),
    .I1(x19_y29),
    .I2(x20_y24),
    .I3(x20_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101010011000)
) lut_23_25 (
    .O(x23_y25),
    .I0(x21_y20),
    .I1(x21_y25),
    .I2(x21_y20),
    .I3(x20_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001011100111)
) lut_24_25 (
    .O(x24_y25),
    .I0(1'b0),
    .I1(x22_y30),
    .I2(x22_y29),
    .I3(x22_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011010100001)
) lut_25_25 (
    .O(x25_y25),
    .I0(x23_y22),
    .I1(x22_y30),
    .I2(x22_y30),
    .I3(x22_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100010100011)
) lut_26_25 (
    .O(x26_y25),
    .I0(x23_y20),
    .I1(x23_y29),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100101001001)
) lut_27_25 (
    .O(x27_y25),
    .I0(x25_y24),
    .I1(x24_y22),
    .I2(1'b0),
    .I3(x24_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011001001111)
) lut_28_25 (
    .O(x28_y25),
    .I0(x26_y23),
    .I1(1'b0),
    .I2(x25_y23),
    .I3(x25_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001111001110)
) lut_29_25 (
    .O(x29_y25),
    .I0(x26_y20),
    .I1(x26_y26),
    .I2(x27_y23),
    .I3(x26_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010000010010)
) lut_30_25 (
    .O(x30_y25),
    .I0(x27_y21),
    .I1(x28_y29),
    .I2(1'b0),
    .I3(x27_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100011101101)
) lut_31_25 (
    .O(x31_y25),
    .I0(x28_y29),
    .I1(x28_y30),
    .I2(x28_y24),
    .I3(x28_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111100000011)
) lut_32_25 (
    .O(x32_y25),
    .I0(x29_y28),
    .I1(x30_y22),
    .I2(x30_y29),
    .I3(x30_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011111110111)
) lut_33_25 (
    .O(x33_y25),
    .I0(x30_y25),
    .I1(x30_y26),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010100100110)
) lut_34_25 (
    .O(x34_y25),
    .I0(x32_y20),
    .I1(x32_y26),
    .I2(x31_y28),
    .I3(x32_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001100110001)
) lut_35_25 (
    .O(x35_y25),
    .I0(x33_y25),
    .I1(x33_y21),
    .I2(x32_y25),
    .I3(x32_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100111011111)
) lut_36_25 (
    .O(x36_y25),
    .I0(1'b0),
    .I1(x34_y25),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010111101000)
) lut_37_25 (
    .O(x37_y25),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x35_y20),
    .I3(x35_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010110001110)
) lut_38_25 (
    .O(x38_y25),
    .I0(x35_y24),
    .I1(x36_y28),
    .I2(x35_y26),
    .I3(x35_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000011011000)
) lut_39_25 (
    .O(x39_y25),
    .I0(x37_y29),
    .I1(1'b0),
    .I2(x37_y20),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001010010101)
) lut_40_25 (
    .O(x40_y25),
    .I0(1'b0),
    .I1(x38_y25),
    .I2(1'b0),
    .I3(x37_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101010011111)
) lut_41_25 (
    .O(x41_y25),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x39_y23),
    .I3(x38_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100101110011)
) lut_42_25 (
    .O(x42_y25),
    .I0(x39_y24),
    .I1(x39_y30),
    .I2(x40_y23),
    .I3(x39_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011101111011)
) lut_43_25 (
    .O(x43_y25),
    .I0(x41_y27),
    .I1(1'b0),
    .I2(x41_y20),
    .I3(x41_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001110010001)
) lut_44_25 (
    .O(x44_y25),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x42_y24),
    .I3(x41_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010010100000)
) lut_45_25 (
    .O(x45_y25),
    .I0(x43_y24),
    .I1(x42_y27),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100000111011)
) lut_46_25 (
    .O(x46_y25),
    .I0(x44_y25),
    .I1(1'b0),
    .I2(x43_y28),
    .I3(x44_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001011011011)
) lut_47_25 (
    .O(x47_y25),
    .I0(x45_y30),
    .I1(1'b0),
    .I2(x44_y20),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111011101101)
) lut_48_25 (
    .O(x48_y25),
    .I0(1'b0),
    .I1(x45_y27),
    .I2(x46_y26),
    .I3(x46_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111010110011)
) lut_49_25 (
    .O(x49_y25),
    .I0(x46_y29),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101011011010)
) lut_50_25 (
    .O(x50_y25),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x48_y30),
    .I3(x48_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111010111110)
) lut_51_25 (
    .O(x51_y25),
    .I0(1'b0),
    .I1(x49_y22),
    .I2(x49_y29),
    .I3(x48_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011001110111)
) lut_52_25 (
    .O(x52_y25),
    .I0(x49_y25),
    .I1(x49_y25),
    .I2(x49_y29),
    .I3(x49_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001011111010)
) lut_53_25 (
    .O(x53_y25),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x50_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010000010001)
) lut_54_25 (
    .O(x54_y25),
    .I0(x52_y26),
    .I1(1'b0),
    .I2(x51_y24),
    .I3(x51_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110110111111)
) lut_55_25 (
    .O(x55_y25),
    .I0(1'b0),
    .I1(x52_y20),
    .I2(x52_y29),
    .I3(x53_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110011111000)
) lut_56_25 (
    .O(x56_y25),
    .I0(x53_y28),
    .I1(x54_y28),
    .I2(x53_y26),
    .I3(x53_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011011001000)
) lut_57_25 (
    .O(x57_y25),
    .I0(1'b0),
    .I1(x54_y23),
    .I2(x55_y27),
    .I3(x54_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100011011111)
) lut_58_25 (
    .O(x58_y25),
    .I0(x56_y23),
    .I1(x56_y22),
    .I2(x55_y21),
    .I3(x56_y20)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000110010100)
) lut_59_25 (
    .O(x59_y25),
    .I0(x56_y21),
    .I1(x56_y29),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001010111111)
) lut_60_25 (
    .O(x60_y25),
    .I0(x58_y20),
    .I1(x58_y25),
    .I2(x57_y22),
    .I3(x58_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010001110010)
) lut_61_25 (
    .O(x61_y25),
    .I0(x59_y26),
    .I1(x58_y23),
    .I2(x58_y22),
    .I3(x58_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101011100000)
) lut_62_25 (
    .O(x62_y25),
    .I0(x59_y29),
    .I1(x60_y27),
    .I2(x59_y27),
    .I3(x59_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100110000101)
) lut_0_26 (
    .O(x0_y26),
    .I0(1'b0),
    .I1(in8),
    .I2(1'b0),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100010001010)
) lut_1_26 (
    .O(x1_y26),
    .I0(1'b0),
    .I1(in3),
    .I2(1'b0),
    .I3(in6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000000100110)
) lut_2_26 (
    .O(x2_y26),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100001011101)
) lut_3_26 (
    .O(x3_y26),
    .I0(in8),
    .I1(1'b0),
    .I2(in2),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100010110000)
) lut_4_26 (
    .O(x4_y26),
    .I0(1'b0),
    .I1(x2_y24),
    .I2(x2_y28),
    .I3(x2_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010001000000)
) lut_5_26 (
    .O(x5_y26),
    .I0(x3_y26),
    .I1(x3_y25),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000100000001)
) lut_6_26 (
    .O(x6_y26),
    .I0(x3_y22),
    .I1(x3_y26),
    .I2(x3_y24),
    .I3(x3_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100001010110)
) lut_7_26 (
    .O(x7_y26),
    .I0(1'b0),
    .I1(x5_y24),
    .I2(x5_y23),
    .I3(x4_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001001110010)
) lut_8_26 (
    .O(x8_y26),
    .I0(x6_y29),
    .I1(x5_y24),
    .I2(x5_y29),
    .I3(x5_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011111001010)
) lut_9_26 (
    .O(x9_y26),
    .I0(x7_y26),
    .I1(x7_y24),
    .I2(x5_y29),
    .I3(x5_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000110110100)
) lut_10_26 (
    .O(x10_y26),
    .I0(x7_y30),
    .I1(1'b0),
    .I2(x7_y23),
    .I3(x7_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110100001011)
) lut_11_26 (
    .O(x11_y26),
    .I0(x8_y23),
    .I1(1'b0),
    .I2(x8_y29),
    .I3(x8_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000110000100)
) lut_12_26 (
    .O(x12_y26),
    .I0(x9_y25),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x9_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101111110100)
) lut_13_26 (
    .O(x13_y26),
    .I0(x10_y25),
    .I1(x11_y28),
    .I2(x10_y22),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110010101000)
) lut_14_26 (
    .O(x14_y26),
    .I0(1'b0),
    .I1(x11_y26),
    .I2(x12_y23),
    .I3(x11_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101110110010)
) lut_15_26 (
    .O(x15_y26),
    .I0(x12_y29),
    .I1(x12_y29),
    .I2(x13_y25),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111011110111)
) lut_16_26 (
    .O(x16_y26),
    .I0(x13_y23),
    .I1(x13_y29),
    .I2(x14_y26),
    .I3(x14_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111110010110)
) lut_17_26 (
    .O(x17_y26),
    .I0(1'b0),
    .I1(x15_y21),
    .I2(x14_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111101111111)
) lut_18_26 (
    .O(x18_y26),
    .I0(x16_y24),
    .I1(x16_y29),
    .I2(x15_y29),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110001101101)
) lut_19_26 (
    .O(x19_y26),
    .I0(x16_y30),
    .I1(x16_y22),
    .I2(1'b0),
    .I3(x17_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000111110101)
) lut_20_26 (
    .O(x20_y26),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x17_y27),
    .I3(x18_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111101011000)
) lut_21_26 (
    .O(x21_y26),
    .I0(x18_y27),
    .I1(x19_y30),
    .I2(x18_y24),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101111111000)
) lut_22_26 (
    .O(x22_y26),
    .I0(x20_y28),
    .I1(x20_y24),
    .I2(1'b0),
    .I3(x19_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001011001100)
) lut_23_26 (
    .O(x23_y26),
    .I0(x21_y30),
    .I1(1'b0),
    .I2(x21_y25),
    .I3(x21_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001110000101)
) lut_24_26 (
    .O(x24_y26),
    .I0(x21_y27),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x22_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100011100110)
) lut_25_26 (
    .O(x25_y26),
    .I0(x23_y21),
    .I1(x23_y30),
    .I2(x22_y21),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100101110010)
) lut_26_26 (
    .O(x26_y26),
    .I0(x23_y24),
    .I1(1'b0),
    .I2(x24_y23),
    .I3(x23_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100000110011)
) lut_27_26 (
    .O(x27_y26),
    .I0(x24_y28),
    .I1(1'b0),
    .I2(x24_y28),
    .I3(x25_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011100001110)
) lut_28_26 (
    .O(x28_y26),
    .I0(x26_y22),
    .I1(x25_y31),
    .I2(x25_y29),
    .I3(x26_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110100000011)
) lut_29_26 (
    .O(x29_y26),
    .I0(x27_y24),
    .I1(x27_y31),
    .I2(x27_y23),
    .I3(x27_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100111110100)
) lut_30_26 (
    .O(x30_y26),
    .I0(x28_y23),
    .I1(x27_y23),
    .I2(x27_y21),
    .I3(x28_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001000000001)
) lut_31_26 (
    .O(x31_y26),
    .I0(1'b0),
    .I1(x29_y22),
    .I2(1'b0),
    .I3(x28_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011010001101)
) lut_32_26 (
    .O(x32_y26),
    .I0(x30_y31),
    .I1(x29_y23),
    .I2(1'b0),
    .I3(x29_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000101010100)
) lut_33_26 (
    .O(x33_y26),
    .I0(x31_y26),
    .I1(x31_y29),
    .I2(x30_y24),
    .I3(x30_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011110001010)
) lut_34_26 (
    .O(x34_y26),
    .I0(x32_y26),
    .I1(x32_y26),
    .I2(x31_y26),
    .I3(x32_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110011100101)
) lut_35_26 (
    .O(x35_y26),
    .I0(x33_y24),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x33_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010010101111)
) lut_36_26 (
    .O(x36_y26),
    .I0(x34_y23),
    .I1(x33_y25),
    .I2(x33_y21),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101110101100)
) lut_37_26 (
    .O(x37_y26),
    .I0(1'b0),
    .I1(x35_y29),
    .I2(x34_y25),
    .I3(x35_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110101011110)
) lut_38_26 (
    .O(x38_y26),
    .I0(x36_y27),
    .I1(x35_y27),
    .I2(x35_y25),
    .I3(x36_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011111010000)
) lut_39_26 (
    .O(x39_y26),
    .I0(x36_y27),
    .I1(1'b0),
    .I2(x37_y23),
    .I3(x36_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100000100101)
) lut_40_26 (
    .O(x40_y26),
    .I0(x38_y29),
    .I1(x38_y28),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000101010001)
) lut_41_26 (
    .O(x41_y26),
    .I0(1'b0),
    .I1(x39_y22),
    .I2(x38_y23),
    .I3(x38_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011111010000)
) lut_42_26 (
    .O(x42_y26),
    .I0(x40_y26),
    .I1(1'b0),
    .I2(x39_y23),
    .I3(x40_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000000111011)
) lut_43_26 (
    .O(x43_y26),
    .I0(x40_y28),
    .I1(x40_y28),
    .I2(x40_y28),
    .I3(x40_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010011110001)
) lut_44_26 (
    .O(x44_y26),
    .I0(x42_y30),
    .I1(x41_y28),
    .I2(x41_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011001100001)
) lut_45_26 (
    .O(x45_y26),
    .I0(x43_y23),
    .I1(x43_y26),
    .I2(x42_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000110010000)
) lut_46_26 (
    .O(x46_y26),
    .I0(1'b0),
    .I1(x44_y27),
    .I2(x44_y22),
    .I3(x44_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001100101011)
) lut_47_26 (
    .O(x47_y26),
    .I0(x44_y23),
    .I1(x45_y24),
    .I2(x45_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100111010100)
) lut_48_26 (
    .O(x48_y26),
    .I0(x45_y22),
    .I1(x45_y28),
    .I2(x46_y22),
    .I3(x45_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010011100011)
) lut_49_26 (
    .O(x49_y26),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x47_y25),
    .I3(x47_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100100001110)
) lut_50_26 (
    .O(x50_y26),
    .I0(x47_y24),
    .I1(x47_y24),
    .I2(x48_y31),
    .I3(x47_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111110101100)
) lut_51_26 (
    .O(x51_y26),
    .I0(x49_y24),
    .I1(x48_y26),
    .I2(x49_y28),
    .I3(x49_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101110000010)
) lut_52_26 (
    .O(x52_y26),
    .I0(x49_y29),
    .I1(x50_y31),
    .I2(x50_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100100000010)
) lut_53_26 (
    .O(x53_y26),
    .I0(x51_y23),
    .I1(x50_y30),
    .I2(x51_y30),
    .I3(x50_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110101000111)
) lut_54_26 (
    .O(x54_y26),
    .I0(x51_y23),
    .I1(x51_y26),
    .I2(x51_y28),
    .I3(x51_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011100000001)
) lut_55_26 (
    .O(x55_y26),
    .I0(x53_y24),
    .I1(1'b0),
    .I2(x52_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001001000100)
) lut_56_26 (
    .O(x56_y26),
    .I0(x54_y27),
    .I1(x53_y22),
    .I2(1'b0),
    .I3(x53_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001010001000)
) lut_57_26 (
    .O(x57_y26),
    .I0(x55_y21),
    .I1(x54_y26),
    .I2(x55_y29),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110111001110)
) lut_58_26 (
    .O(x58_y26),
    .I0(x56_y23),
    .I1(x55_y25),
    .I2(x56_y24),
    .I3(x56_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011011000100)
) lut_59_26 (
    .O(x59_y26),
    .I0(x56_y24),
    .I1(1'b0),
    .I2(x56_y22),
    .I3(x56_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100100100011)
) lut_60_26 (
    .O(x60_y26),
    .I0(1'b0),
    .I1(x57_y28),
    .I2(x58_y21),
    .I3(x58_y21)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001110001011)
) lut_61_26 (
    .O(x61_y26),
    .I0(x58_y22),
    .I1(x58_y29),
    .I2(x58_y21),
    .I3(x59_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110110000010)
) lut_62_26 (
    .O(x62_y26),
    .I0(x59_y24),
    .I1(x59_y26),
    .I2(1'b0),
    .I3(x60_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001110000000)
) lut_0_27 (
    .O(x0_y27),
    .I0(in9),
    .I1(1'b0),
    .I2(in7),
    .I3(in9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010111101010)
) lut_1_27 (
    .O(x1_y27),
    .I0(1'b0),
    .I1(in9),
    .I2(in6),
    .I3(in9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110100001110)
) lut_2_27 (
    .O(x2_y27),
    .I0(in4),
    .I1(in9),
    .I2(in9),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001010010010)
) lut_3_27 (
    .O(x3_y27),
    .I0(x1_y28),
    .I1(x1_y31),
    .I2(in3),
    .I3(in7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101001011010)
) lut_4_27 (
    .O(x4_y27),
    .I0(x1_y22),
    .I1(x1_y24),
    .I2(x1_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111101101010)
) lut_5_27 (
    .O(x5_y27),
    .I0(x2_y25),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100110110110)
) lut_6_27 (
    .O(x6_y27),
    .I0(x3_y26),
    .I1(x3_y25),
    .I2(1'b0),
    .I3(x4_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001101000000)
) lut_7_27 (
    .O(x7_y27),
    .I0(x4_y32),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x5_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101011100000)
) lut_8_27 (
    .O(x8_y27),
    .I0(x5_y27),
    .I1(x5_y31),
    .I2(x6_y27),
    .I3(x6_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101011001011)
) lut_9_27 (
    .O(x9_y27),
    .I0(x7_y30),
    .I1(x6_y27),
    .I2(x6_y27),
    .I3(x6_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000001011100)
) lut_10_27 (
    .O(x10_y27),
    .I0(x8_y31),
    .I1(x7_y22),
    .I2(x8_y24),
    .I3(x7_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110011111001)
) lut_11_27 (
    .O(x11_y27),
    .I0(x9_y30),
    .I1(x8_y25),
    .I2(x8_y26),
    .I3(x8_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011110101100)
) lut_12_27 (
    .O(x12_y27),
    .I0(1'b0),
    .I1(x9_y32),
    .I2(x9_y29),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011100110101)
) lut_13_27 (
    .O(x13_y27),
    .I0(1'b0),
    .I1(x11_y22),
    .I2(1'b0),
    .I3(x10_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110110110111)
) lut_14_27 (
    .O(x14_y27),
    .I0(x11_y23),
    .I1(x11_y26),
    .I2(x11_y29),
    .I3(x12_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000001101011)
) lut_15_27 (
    .O(x15_y27),
    .I0(x13_y32),
    .I1(x12_y32),
    .I2(1'b0),
    .I3(x13_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010001001000)
) lut_16_27 (
    .O(x16_y27),
    .I0(x13_y29),
    .I1(x14_y27),
    .I2(x13_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010100101011)
) lut_17_27 (
    .O(x17_y27),
    .I0(x15_y27),
    .I1(1'b0),
    .I2(x15_y25),
    .I3(x14_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011110011111)
) lut_18_27 (
    .O(x18_y27),
    .I0(x16_y32),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011010101001)
) lut_19_27 (
    .O(x19_y27),
    .I0(1'b0),
    .I1(x16_y32),
    .I2(x16_y27),
    .I3(x17_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000100111001)
) lut_20_27 (
    .O(x20_y27),
    .I0(x17_y24),
    .I1(x17_y29),
    .I2(x17_y25),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010011000101)
) lut_21_27 (
    .O(x21_y27),
    .I0(x19_y30),
    .I1(x18_y29),
    .I2(1'b0),
    .I3(x18_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110100010111)
) lut_22_27 (
    .O(x22_y27),
    .I0(x20_y30),
    .I1(x20_y26),
    .I2(x19_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000101000000)
) lut_23_27 (
    .O(x23_y27),
    .I0(x20_y29),
    .I1(x20_y27),
    .I2(1'b0),
    .I3(x21_y22)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010000110001)
) lut_24_27 (
    .O(x24_y27),
    .I0(1'b0),
    .I1(x22_y27),
    .I2(x22_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000010100101)
) lut_25_27 (
    .O(x25_y27),
    .I0(x23_y28),
    .I1(x23_y26),
    .I2(1'b0),
    .I3(x23_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001111101101)
) lut_26_27 (
    .O(x26_y27),
    .I0(x23_y23),
    .I1(x23_y24),
    .I2(x23_y28),
    .I3(x23_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001011010010)
) lut_27_27 (
    .O(x27_y27),
    .I0(x24_y24),
    .I1(x24_y27),
    .I2(x24_y24),
    .I3(x25_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000010001110)
) lut_28_27 (
    .O(x28_y27),
    .I0(1'b0),
    .I1(x26_y32),
    .I2(x25_y26),
    .I3(x26_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101111011101)
) lut_29_27 (
    .O(x29_y27),
    .I0(x26_y30),
    .I1(1'b0),
    .I2(x27_y31),
    .I3(x27_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011001010001)
) lut_30_27 (
    .O(x30_y27),
    .I0(x27_y28),
    .I1(x27_y30),
    .I2(1'b0),
    .I3(x28_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000010111001)
) lut_31_27 (
    .O(x31_y27),
    .I0(x28_y25),
    .I1(x28_y26),
    .I2(x28_y26),
    .I3(x28_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000010001111)
) lut_32_27 (
    .O(x32_y27),
    .I0(1'b0),
    .I1(x30_y28),
    .I2(x29_y22),
    .I3(x30_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000100001100)
) lut_33_27 (
    .O(x33_y27),
    .I0(x31_y30),
    .I1(1'b0),
    .I2(x31_y22),
    .I3(x31_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011100101101)
) lut_34_27 (
    .O(x34_y27),
    .I0(1'b0),
    .I1(x31_y32),
    .I2(x32_y31),
    .I3(x31_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100100010010)
) lut_35_27 (
    .O(x35_y27),
    .I0(x33_y27),
    .I1(1'b0),
    .I2(x33_y23),
    .I3(x33_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011110111111)
) lut_36_27 (
    .O(x36_y27),
    .I0(1'b0),
    .I1(x34_y24),
    .I2(1'b0),
    .I3(x34_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001100000011)
) lut_37_27 (
    .O(x37_y27),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x35_y29),
    .I3(x35_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111101110010)
) lut_38_27 (
    .O(x38_y27),
    .I0(x35_y26),
    .I1(x35_y24),
    .I2(x36_y31),
    .I3(x35_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111000000010)
) lut_39_27 (
    .O(x39_y27),
    .I0(x37_y22),
    .I1(x36_y28),
    .I2(x37_y23),
    .I3(x37_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110100111011)
) lut_40_27 (
    .O(x40_y27),
    .I0(x37_y24),
    .I1(x37_y24),
    .I2(x38_y28),
    .I3(x38_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011101001010)
) lut_41_27 (
    .O(x41_y27),
    .I0(x39_y26),
    .I1(x38_y27),
    .I2(x38_y32),
    .I3(x38_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111111000110)
) lut_42_27 (
    .O(x42_y27),
    .I0(x39_y26),
    .I1(1'b0),
    .I2(x40_y22),
    .I3(x39_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110011101101)
) lut_43_27 (
    .O(x43_y27),
    .I0(x41_y27),
    .I1(x40_y23),
    .I2(x41_y26),
    .I3(x41_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011111000110)
) lut_44_27 (
    .O(x44_y27),
    .I0(x41_y24),
    .I1(1'b0),
    .I2(x41_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101100010101)
) lut_45_27 (
    .O(x45_y27),
    .I0(1'b0),
    .I1(x43_y30),
    .I2(x43_y27),
    .I3(x42_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001100010111)
) lut_46_27 (
    .O(x46_y27),
    .I0(x44_y31),
    .I1(x44_y22),
    .I2(x44_y25),
    .I3(x44_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001010011111)
) lut_47_27 (
    .O(x47_y27),
    .I0(x45_y32),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x44_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100010011100)
) lut_48_27 (
    .O(x48_y27),
    .I0(x45_y27),
    .I1(x45_y27),
    .I2(x45_y31),
    .I3(x46_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100111101111)
) lut_49_27 (
    .O(x49_y27),
    .I0(x46_y24),
    .I1(x46_y30),
    .I2(x46_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000100001111)
) lut_50_27 (
    .O(x50_y27),
    .I0(x48_y25),
    .I1(x47_y23),
    .I2(x47_y29),
    .I3(x47_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111010011010)
) lut_51_27 (
    .O(x51_y27),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x48_y25),
    .I3(x49_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000001010101)
) lut_52_27 (
    .O(x52_y27),
    .I0(x50_y32),
    .I1(x49_y23),
    .I2(1'b0),
    .I3(x49_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011101101001)
) lut_53_27 (
    .O(x53_y27),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x51_y29),
    .I3(x50_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110110001000)
) lut_54_27 (
    .O(x54_y27),
    .I0(x52_y31),
    .I1(x52_y25),
    .I2(1'b0),
    .I3(x52_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110101011001)
) lut_55_27 (
    .O(x55_y27),
    .I0(x52_y26),
    .I1(1'b0),
    .I2(x53_y31),
    .I3(x52_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000110111111)
) lut_56_27 (
    .O(x56_y27),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x54_y31),
    .I3(x54_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010011111010)
) lut_57_27 (
    .O(x57_y27),
    .I0(1'b0),
    .I1(x55_y28),
    .I2(1'b0),
    .I3(x55_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000101011010)
) lut_58_27 (
    .O(x58_y27),
    .I0(x56_y25),
    .I1(x55_y31),
    .I2(1'b0),
    .I3(x56_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001000000111)
) lut_59_27 (
    .O(x59_y27),
    .I0(x56_y30),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x57_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000010101100)
) lut_60_27 (
    .O(x60_y27),
    .I0(x57_y29),
    .I1(x57_y30),
    .I2(x57_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011111110111)
) lut_61_27 (
    .O(x61_y27),
    .I0(x58_y27),
    .I1(x59_y22),
    .I2(x59_y25),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011001011110)
) lut_62_27 (
    .O(x62_y27),
    .I0(x60_y23),
    .I1(x60_y29),
    .I2(x60_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100001000100)
) lut_0_28 (
    .O(x0_y28),
    .I0(in8),
    .I1(in3),
    .I2(in3),
    .I3(in5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111101001111)
) lut_1_28 (
    .O(x1_y28),
    .I0(in3),
    .I1(in6),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110011110110)
) lut_2_28 (
    .O(x2_y28),
    .I0(in9),
    .I1(in9),
    .I2(in6),
    .I3(in7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010100001001)
) lut_3_28 (
    .O(x3_y28),
    .I0(x1_y25),
    .I1(x1_y24),
    .I2(x1_y23),
    .I3(x1_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110010000010)
) lut_4_28 (
    .O(x4_y28),
    .I0(x1_y31),
    .I1(x2_y32),
    .I2(x1_y25),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100011110110)
) lut_5_28 (
    .O(x5_y28),
    .I0(x3_y24),
    .I1(x3_y32),
    .I2(x3_y28),
    .I3(x3_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000011001111)
) lut_6_28 (
    .O(x6_y28),
    .I0(x3_y33),
    .I1(x4_y27),
    .I2(x3_y26),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110000110101)
) lut_7_28 (
    .O(x7_y28),
    .I0(x5_y31),
    .I1(x5_y27),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001000101000)
) lut_8_28 (
    .O(x8_y28),
    .I0(x6_y32),
    .I1(x5_y26),
    .I2(x5_y24),
    .I3(x5_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111000101001)
) lut_9_28 (
    .O(x9_y28),
    .I0(x6_y31),
    .I1(x6_y29),
    .I2(x5_y24),
    .I3(x5_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111101011101)
) lut_10_28 (
    .O(x10_y28),
    .I0(x8_y33),
    .I1(1'b0),
    .I2(x8_y31),
    .I3(x7_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101000001010)
) lut_11_28 (
    .O(x11_y28),
    .I0(x9_y32),
    .I1(x8_y28),
    .I2(1'b0),
    .I3(x8_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101011101111)
) lut_12_28 (
    .O(x12_y28),
    .I0(1'b0),
    .I1(x10_y27),
    .I2(x9_y28),
    .I3(x10_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011000001011)
) lut_13_28 (
    .O(x13_y28),
    .I0(x10_y23),
    .I1(1'b0),
    .I2(x11_y29),
    .I3(x10_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100001001000)
) lut_14_28 (
    .O(x14_y28),
    .I0(x11_y31),
    .I1(1'b0),
    .I2(x11_y23),
    .I3(x11_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011010010110)
) lut_15_28 (
    .O(x15_y28),
    .I0(x13_y27),
    .I1(x13_y31),
    .I2(x12_y30),
    .I3(x12_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110100111100)
) lut_16_28 (
    .O(x16_y28),
    .I0(x14_y32),
    .I1(x14_y30),
    .I2(x13_y27),
    .I3(x14_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011111010010)
) lut_17_28 (
    .O(x17_y28),
    .I0(x14_y27),
    .I1(x14_y30),
    .I2(x14_y28),
    .I3(x14_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101001110111)
) lut_18_28 (
    .O(x18_y28),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x15_y26),
    .I3(x16_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100000100110)
) lut_19_28 (
    .O(x19_y28),
    .I0(1'b0),
    .I1(x16_y27),
    .I2(1'b0),
    .I3(x17_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110111100010)
) lut_20_28 (
    .O(x20_y28),
    .I0(1'b0),
    .I1(x17_y25),
    .I2(x17_y27),
    .I3(x18_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010111010010)
) lut_21_28 (
    .O(x21_y28),
    .I0(x19_y27),
    .I1(1'b0),
    .I2(x19_y30),
    .I3(x19_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010000111000)
) lut_22_28 (
    .O(x22_y28),
    .I0(x19_y32),
    .I1(1'b0),
    .I2(x19_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010011111110)
) lut_23_28 (
    .O(x23_y28),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x20_y27),
    .I3(x21_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111100110100)
) lut_24_28 (
    .O(x24_y28),
    .I0(x22_y30),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111010110111)
) lut_25_28 (
    .O(x25_y28),
    .I0(x23_y23),
    .I1(x23_y23),
    .I2(x23_y29),
    .I3(x23_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100111111010)
) lut_26_28 (
    .O(x26_y28),
    .I0(x23_y32),
    .I1(x23_y26),
    .I2(1'b0),
    .I3(x23_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010100101100)
) lut_27_28 (
    .O(x27_y28),
    .I0(x24_y29),
    .I1(x25_y23),
    .I2(1'b0),
    .I3(x24_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000011010110)
) lut_28_28 (
    .O(x28_y28),
    .I0(x25_y23),
    .I1(x25_y24),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010111001110)
) lut_29_28 (
    .O(x29_y28),
    .I0(1'b0),
    .I1(x26_y32),
    .I2(x27_y23),
    .I3(x27_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010100010111)
) lut_30_28 (
    .O(x30_y28),
    .I0(x27_y31),
    .I1(x27_y27),
    .I2(x27_y28),
    .I3(x28_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010110010111)
) lut_31_28 (
    .O(x31_y28),
    .I0(x29_y23),
    .I1(x29_y25),
    .I2(x28_y31),
    .I3(x28_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100100101011)
) lut_32_28 (
    .O(x32_y28),
    .I0(x29_y24),
    .I1(x29_y31),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011111110111)
) lut_33_28 (
    .O(x33_y28),
    .I0(x31_y27),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x31_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110111111111)
) lut_34_28 (
    .O(x34_y28),
    .I0(x32_y30),
    .I1(x31_y31),
    .I2(x32_y33),
    .I3(x32_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011111111001)
) lut_35_28 (
    .O(x35_y28),
    .I0(x32_y25),
    .I1(x32_y24),
    .I2(x32_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101111101010)
) lut_36_28 (
    .O(x36_y28),
    .I0(x34_y26),
    .I1(1'b0),
    .I2(x33_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110101011000)
) lut_37_28 (
    .O(x37_y28),
    .I0(x35_y29),
    .I1(x34_y28),
    .I2(1'b0),
    .I3(x34_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011101000000)
) lut_38_28 (
    .O(x38_y28),
    .I0(x35_y26),
    .I1(1'b0),
    .I2(x35_y23),
    .I3(x36_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011001001101)
) lut_39_28 (
    .O(x39_y28),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111101011111)
) lut_40_28 (
    .O(x40_y28),
    .I0(x38_y26),
    .I1(x38_y25),
    .I2(x38_y24),
    .I3(x38_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010100000110)
) lut_41_28 (
    .O(x41_y28),
    .I0(x38_y32),
    .I1(x38_y28),
    .I2(x39_y30),
    .I3(x38_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110101110111)
) lut_42_28 (
    .O(x42_y28),
    .I0(x40_y32),
    .I1(x39_y32),
    .I2(x40_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011000010011)
) lut_43_28 (
    .O(x43_y28),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x41_y30),
    .I3(x40_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001000011110)
) lut_44_28 (
    .O(x44_y28),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x41_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110001100101)
) lut_45_28 (
    .O(x45_y28),
    .I0(1'b0),
    .I1(x42_y23),
    .I2(x43_y28),
    .I3(x42_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100101011001)
) lut_46_28 (
    .O(x46_y28),
    .I0(x44_y25),
    .I1(x44_y31),
    .I2(x43_y32),
    .I3(x44_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110101101110)
) lut_47_28 (
    .O(x47_y28),
    .I0(1'b0),
    .I1(x44_y24),
    .I2(x44_y29),
    .I3(x44_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001101011101)
) lut_48_28 (
    .O(x48_y28),
    .I0(1'b0),
    .I1(x46_y29),
    .I2(1'b0),
    .I3(x45_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100010010010)
) lut_49_28 (
    .O(x49_y28),
    .I0(1'b0),
    .I1(x46_y26),
    .I2(1'b0),
    .I3(x47_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110110011000)
) lut_50_28 (
    .O(x50_y28),
    .I0(x48_y29),
    .I1(x47_y25),
    .I2(x48_y23),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101100010100)
) lut_51_28 (
    .O(x51_y28),
    .I0(x48_y31),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010000111010)
) lut_52_28 (
    .O(x52_y28),
    .I0(x49_y33),
    .I1(x49_y24),
    .I2(x49_y28),
    .I3(x49_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001010011111)
) lut_53_28 (
    .O(x53_y28),
    .I0(x50_y26),
    .I1(x51_y23),
    .I2(x50_y26),
    .I3(x51_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111011100010)
) lut_54_28 (
    .O(x54_y28),
    .I0(x52_y29),
    .I1(x52_y27),
    .I2(x51_y24),
    .I3(x51_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101110000100)
) lut_55_28 (
    .O(x55_y28),
    .I0(x53_y30),
    .I1(x53_y26),
    .I2(x52_y27),
    .I3(x52_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111000110111)
) lut_56_28 (
    .O(x56_y28),
    .I0(x53_y29),
    .I1(x54_y24),
    .I2(x53_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110110111101)
) lut_57_28 (
    .O(x57_y28),
    .I0(x54_y31),
    .I1(x55_y30),
    .I2(x54_y25),
    .I3(x54_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010100000100)
) lut_58_28 (
    .O(x58_y28),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x55_y31),
    .I3(x55_y23)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100110110010)
) lut_59_28 (
    .O(x59_y28),
    .I0(x56_y25),
    .I1(x57_y31),
    .I2(1'b0),
    .I3(x56_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101010101010)
) lut_60_28 (
    .O(x60_y28),
    .I0(1'b0),
    .I1(x57_y23),
    .I2(x57_y32),
    .I3(x57_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101110001000)
) lut_61_28 (
    .O(x61_y28),
    .I0(x58_y25),
    .I1(x59_y28),
    .I2(x58_y33),
    .I3(x59_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010011101000)
) lut_62_28 (
    .O(x62_y28),
    .I0(x59_y26),
    .I1(x60_y29),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100000110000)
) lut_0_29 (
    .O(x0_y29),
    .I0(1'b0),
    .I1(in5),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110100001111)
) lut_1_29 (
    .O(x1_y29),
    .I0(in6),
    .I1(in4),
    .I2(in2),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001101001110)
) lut_2_29 (
    .O(x2_y29),
    .I0(in3),
    .I1(in4),
    .I2(in8),
    .I3(in7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100100110010)
) lut_3_29 (
    .O(x3_y29),
    .I0(in1),
    .I1(1'b0),
    .I2(in4),
    .I3(x1_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100010110111)
) lut_4_29 (
    .O(x4_y29),
    .I0(x2_y34),
    .I1(x1_y26),
    .I2(x1_y24),
    .I3(x2_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000000100110)
) lut_5_29 (
    .O(x5_y29),
    .I0(x3_y28),
    .I1(x3_y29),
    .I2(x3_y27),
    .I3(x2_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100011010110)
) lut_6_29 (
    .O(x6_y29),
    .I0(x4_y26),
    .I1(x4_y31),
    .I2(x4_y28),
    .I3(x3_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010110110000)
) lut_7_29 (
    .O(x7_y29),
    .I0(x5_y34),
    .I1(x5_y27),
    .I2(x5_y34),
    .I3(x5_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001100101000)
) lut_8_29 (
    .O(x8_y29),
    .I0(x5_y33),
    .I1(x5_y28),
    .I2(1'b0),
    .I3(x6_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111101000111)
) lut_9_29 (
    .O(x9_y29),
    .I0(x6_y27),
    .I1(x6_y28),
    .I2(1'b0),
    .I3(x6_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000101000111)
) lut_10_29 (
    .O(x10_y29),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x8_y26),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011011010000)
) lut_11_29 (
    .O(x11_y29),
    .I0(x9_y28),
    .I1(x8_y25),
    .I2(x8_y34),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000110111100)
) lut_12_29 (
    .O(x12_y29),
    .I0(x10_y24),
    .I1(x10_y32),
    .I2(x9_y28),
    .I3(x10_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111101110100)
) lut_13_29 (
    .O(x13_y29),
    .I0(x11_y26),
    .I1(x11_y34),
    .I2(x10_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111000111110)
) lut_14_29 (
    .O(x14_y29),
    .I0(x12_y33),
    .I1(x11_y33),
    .I2(x12_y24),
    .I3(x12_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111000011101)
) lut_15_29 (
    .O(x15_y29),
    .I0(x12_y31),
    .I1(x13_y34),
    .I2(x13_y34),
    .I3(x13_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000111010101)
) lut_16_29 (
    .O(x16_y29),
    .I0(x14_y33),
    .I1(1'b0),
    .I2(x13_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010101010011)
) lut_17_29 (
    .O(x17_y29),
    .I0(x15_y29),
    .I1(x15_y25),
    .I2(x14_y25),
    .I3(x15_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100100010000)
) lut_18_29 (
    .O(x18_y29),
    .I0(x16_y34),
    .I1(x16_y27),
    .I2(x15_y28),
    .I3(x16_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000110001010)
) lut_19_29 (
    .O(x19_y29),
    .I0(1'b0),
    .I1(x16_y34),
    .I2(1'b0),
    .I3(x17_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001100001111)
) lut_20_29 (
    .O(x20_y29),
    .I0(x18_y33),
    .I1(x17_y29),
    .I2(x18_y26),
    .I3(x18_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000001010010)
) lut_21_29 (
    .O(x21_y29),
    .I0(x19_y34),
    .I1(x18_y32),
    .I2(x19_y29),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011001101010)
) lut_22_29 (
    .O(x22_y29),
    .I0(x19_y30),
    .I1(x20_y28),
    .I2(1'b0),
    .I3(x20_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001101010001)
) lut_23_29 (
    .O(x23_y29),
    .I0(x21_y30),
    .I1(x21_y34),
    .I2(x21_y25),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011000100001)
) lut_24_29 (
    .O(x24_y29),
    .I0(x21_y32),
    .I1(x22_y26),
    .I2(x21_y28),
    .I3(x22_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010111110000)
) lut_25_29 (
    .O(x25_y29),
    .I0(x22_y25),
    .I1(x23_y34),
    .I2(x22_y33),
    .I3(x23_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011100100010)
) lut_26_29 (
    .O(x26_y29),
    .I0(x23_y33),
    .I1(x24_y24),
    .I2(x24_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100000001110)
) lut_27_29 (
    .O(x27_y29),
    .I0(x24_y24),
    .I1(1'b0),
    .I2(x25_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011000110001)
) lut_28_29 (
    .O(x28_y29),
    .I0(x26_y25),
    .I1(x25_y27),
    .I2(1'b0),
    .I3(x26_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011011001001)
) lut_29_29 (
    .O(x29_y29),
    .I0(1'b0),
    .I1(x27_y31),
    .I2(1'b0),
    .I3(x27_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101010111111)
) lut_30_29 (
    .O(x30_y29),
    .I0(x28_y27),
    .I1(x27_y24),
    .I2(1'b0),
    .I3(x28_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011010100001)
) lut_31_29 (
    .O(x31_y29),
    .I0(x28_y25),
    .I1(1'b0),
    .I2(x29_y29),
    .I3(x28_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001111111111)
) lut_32_29 (
    .O(x32_y29),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x29_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100111011111)
) lut_33_29 (
    .O(x33_y29),
    .I0(x30_y31),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x31_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011100010011)
) lut_34_29 (
    .O(x34_y29),
    .I0(x31_y24),
    .I1(x31_y31),
    .I2(x31_y31),
    .I3(x32_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111010101101)
) lut_35_29 (
    .O(x35_y29),
    .I0(x33_y28),
    .I1(x33_y26),
    .I2(x33_y33),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100000011111)
) lut_36_29 (
    .O(x36_y29),
    .I0(x33_y28),
    .I1(x34_y28),
    .I2(x33_y25),
    .I3(x33_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011001011100)
) lut_37_29 (
    .O(x37_y29),
    .I0(1'b0),
    .I1(x34_y24),
    .I2(x35_y28),
    .I3(x34_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111101111011)
) lut_38_29 (
    .O(x38_y29),
    .I0(x35_y27),
    .I1(1'b0),
    .I2(x36_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111011011101)
) lut_39_29 (
    .O(x39_y29),
    .I0(x37_y34),
    .I1(x36_y30),
    .I2(x36_y24),
    .I3(x37_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001100101111)
) lut_40_29 (
    .O(x40_y29),
    .I0(x37_y27),
    .I1(x38_y31),
    .I2(1'b0),
    .I3(x37_y24)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100000111101)
) lut_41_29 (
    .O(x41_y29),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x39_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010000001100)
) lut_42_29 (
    .O(x42_y29),
    .I0(x39_y24),
    .I1(1'b0),
    .I2(x39_y34),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010100110011)
) lut_43_29 (
    .O(x43_y29),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x40_y27),
    .I3(x40_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001101011101)
) lut_44_29 (
    .O(x44_y29),
    .I0(x42_y30),
    .I1(x41_y28),
    .I2(x41_y28),
    .I3(x42_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101000011111)
) lut_45_29 (
    .O(x45_y29),
    .I0(x42_y31),
    .I1(x43_y34),
    .I2(x42_y33),
    .I3(x42_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111011010110)
) lut_46_29 (
    .O(x46_y29),
    .I0(x44_y28),
    .I1(x44_y33),
    .I2(x43_y29),
    .I3(x43_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000100100010)
) lut_47_29 (
    .O(x47_y29),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x45_y25),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110110101010)
) lut_48_29 (
    .O(x48_y29),
    .I0(x45_y28),
    .I1(x46_y28),
    .I2(1'b0),
    .I3(x46_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101001101110)
) lut_49_29 (
    .O(x49_y29),
    .I0(x47_y24),
    .I1(x46_y24),
    .I2(1'b0),
    .I3(x47_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011110101011)
) lut_50_29 (
    .O(x50_y29),
    .I0(1'b0),
    .I1(x48_y29),
    .I2(x47_y34),
    .I3(x48_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101000010000)
) lut_51_29 (
    .O(x51_y29),
    .I0(x49_y25),
    .I1(1'b0),
    .I2(x49_y24),
    .I3(x48_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111011101000)
) lut_52_29 (
    .O(x52_y29),
    .I0(x49_y26),
    .I1(x50_y32),
    .I2(x49_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011111001011)
) lut_53_29 (
    .O(x53_y29),
    .I0(x51_y30),
    .I1(x51_y26),
    .I2(x50_y33),
    .I3(x51_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010001000001)
) lut_54_29 (
    .O(x54_y29),
    .I0(x51_y34),
    .I1(x52_y27),
    .I2(x52_y34),
    .I3(x51_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011000101111)
) lut_55_29 (
    .O(x55_y29),
    .I0(x53_y34),
    .I1(x52_y30),
    .I2(x53_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100100111011)
) lut_56_29 (
    .O(x56_y29),
    .I0(1'b0),
    .I1(x53_y33),
    .I2(x54_y26),
    .I3(x54_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100000100101)
) lut_57_29 (
    .O(x57_y29),
    .I0(x54_y34),
    .I1(1'b0),
    .I2(x55_y28),
    .I3(x55_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111111011111)
) lut_58_29 (
    .O(x58_y29),
    .I0(x55_y28),
    .I1(x56_y27),
    .I2(x55_y34),
    .I3(x56_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011101001110)
) lut_59_29 (
    .O(x59_y29),
    .I0(x57_y27),
    .I1(1'b0),
    .I2(x57_y25),
    .I3(x57_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011010101001)
) lut_60_29 (
    .O(x60_y29),
    .I0(x58_y30),
    .I1(x58_y24),
    .I2(x58_y33),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011110100010)
) lut_61_29 (
    .O(x61_y29),
    .I0(x59_y31),
    .I1(1'b0),
    .I2(x58_y27),
    .I3(x59_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111100100111)
) lut_62_29 (
    .O(x62_y29),
    .I0(1'b0),
    .I1(x59_y32),
    .I2(x60_y29),
    .I3(x60_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011010000100)
) lut_0_30 (
    .O(x0_y30),
    .I0(in5),
    .I1(in2),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011101111100)
) lut_1_30 (
    .O(x1_y30),
    .I0(in9),
    .I1(in5),
    .I2(in4),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110101101101)
) lut_2_30 (
    .O(x2_y30),
    .I0(in5),
    .I1(in4),
    .I2(in9),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001111001000)
) lut_3_30 (
    .O(x3_y30),
    .I0(1'b0),
    .I1(x1_y31),
    .I2(1'b0),
    .I3(in6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011101111101)
) lut_4_30 (
    .O(x4_y30),
    .I0(x1_y33),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x1_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011011001011)
) lut_5_30 (
    .O(x5_y30),
    .I0(x3_y25),
    .I1(x3_y26),
    .I2(x3_y33),
    .I3(x2_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110010111001)
) lut_6_30 (
    .O(x6_y30),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x4_y35),
    .I3(x4_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100001000010)
) lut_7_30 (
    .O(x7_y30),
    .I0(x4_y26),
    .I1(1'b0),
    .I2(x4_y35),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000001010011)
) lut_8_30 (
    .O(x8_y30),
    .I0(x5_y31),
    .I1(x6_y34),
    .I2(x6_y33),
    .I3(x5_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110100110101)
) lut_9_30 (
    .O(x9_y30),
    .I0(x7_y29),
    .I1(x7_y31),
    .I2(x6_y33),
    .I3(x5_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101011000011)
) lut_10_30 (
    .O(x10_y30),
    .I0(1'b0),
    .I1(x8_y31),
    .I2(1'b0),
    .I3(x8_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111010110010)
) lut_11_30 (
    .O(x11_y30),
    .I0(x9_y26),
    .I1(1'b0),
    .I2(x8_y25),
    .I3(x8_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111101011111)
) lut_12_30 (
    .O(x12_y30),
    .I0(1'b0),
    .I1(x9_y30),
    .I2(x10_y28),
    .I3(x9_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011001111100)
) lut_13_30 (
    .O(x13_y30),
    .I0(x11_y26),
    .I1(x11_y33),
    .I2(x10_y30),
    .I3(x11_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000110001011)
) lut_14_30 (
    .O(x14_y30),
    .I0(x11_y27),
    .I1(1'b0),
    .I2(x11_y27),
    .I3(x12_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111011000100)
) lut_15_30 (
    .O(x15_y30),
    .I0(1'b0),
    .I1(x13_y26),
    .I2(x12_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111010010111)
) lut_16_30 (
    .O(x16_y30),
    .I0(1'b0),
    .I1(x13_y33),
    .I2(x14_y32),
    .I3(x13_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001101001001)
) lut_17_30 (
    .O(x17_y30),
    .I0(x14_y35),
    .I1(x15_y27),
    .I2(x15_y28),
    .I3(x14_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001100111001)
) lut_18_30 (
    .O(x18_y30),
    .I0(x15_y26),
    .I1(1'b0),
    .I2(x15_y26),
    .I3(x16_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011110110001)
) lut_19_30 (
    .O(x19_y30),
    .I0(x17_y25),
    .I1(x17_y31),
    .I2(x17_y35),
    .I3(x17_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011011011000)
) lut_20_30 (
    .O(x20_y30),
    .I0(x18_y30),
    .I1(1'b0),
    .I2(x18_y34),
    .I3(x17_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010101011111)
) lut_21_30 (
    .O(x21_y30),
    .I0(x19_y26),
    .I1(x18_y29),
    .I2(x18_y29),
    .I3(x18_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110100000011)
) lut_22_30 (
    .O(x22_y30),
    .I0(x20_y34),
    .I1(x19_y29),
    .I2(1'b0),
    .I3(x20_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000101101111)
) lut_23_30 (
    .O(x23_y30),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x21_y35),
    .I3(x20_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100010001111)
) lut_24_30 (
    .O(x24_y30),
    .I0(x21_y27),
    .I1(x22_y28),
    .I2(x22_y27),
    .I3(x22_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000101011001)
) lut_25_30 (
    .O(x25_y30),
    .I0(x22_y30),
    .I1(x22_y25),
    .I2(x23_y33),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010011100000)
) lut_26_30 (
    .O(x26_y30),
    .I0(x24_y35),
    .I1(x24_y32),
    .I2(x23_y34),
    .I3(x23_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010110110100)
) lut_27_30 (
    .O(x27_y30),
    .I0(x25_y28),
    .I1(1'b0),
    .I2(x24_y32),
    .I3(x24_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011100101111)
) lut_28_30 (
    .O(x28_y30),
    .I0(1'b0),
    .I1(x26_y32),
    .I2(x26_y29),
    .I3(x26_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101110000010)
) lut_29_30 (
    .O(x29_y30),
    .I0(1'b0),
    .I1(x26_y31),
    .I2(x27_y27),
    .I3(x27_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111111001000)
) lut_30_30 (
    .O(x30_y30),
    .I0(x27_y35),
    .I1(1'b0),
    .I2(x27_y35),
    .I3(x27_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001010101101)
) lut_31_30 (
    .O(x31_y30),
    .I0(x29_y27),
    .I1(x29_y33),
    .I2(x29_y30),
    .I3(x29_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101111111001)
) lut_32_30 (
    .O(x32_y30),
    .I0(x29_y33),
    .I1(x29_y26),
    .I2(x30_y32),
    .I3(x30_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011101100111)
) lut_33_30 (
    .O(x33_y30),
    .I0(1'b0),
    .I1(x30_y34),
    .I2(x31_y31),
    .I3(x30_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011000110000)
) lut_34_30 (
    .O(x34_y30),
    .I0(1'b0),
    .I1(x31_y27),
    .I2(x31_y31),
    .I3(x31_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000100111000)
) lut_35_30 (
    .O(x35_y30),
    .I0(x33_y28),
    .I1(x32_y29),
    .I2(x33_y30),
    .I3(x33_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011001111110)
) lut_36_30 (
    .O(x36_y30),
    .I0(1'b0),
    .I1(x33_y35),
    .I2(x33_y32),
    .I3(x33_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100000100011)
) lut_37_30 (
    .O(x37_y30),
    .I0(x34_y30),
    .I1(x35_y35),
    .I2(x35_y28),
    .I3(x35_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100101010110)
) lut_38_30 (
    .O(x38_y30),
    .I0(x36_y29),
    .I1(x35_y29),
    .I2(x36_y33),
    .I3(x36_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010010101001)
) lut_39_30 (
    .O(x39_y30),
    .I0(1'b0),
    .I1(x37_y25),
    .I2(x37_y30),
    .I3(x37_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011111011010)
) lut_40_30 (
    .O(x40_y30),
    .I0(x38_y26),
    .I1(x38_y26),
    .I2(x37_y33),
    .I3(x38_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110111011001)
) lut_41_30 (
    .O(x41_y30),
    .I0(x39_y35),
    .I1(x38_y32),
    .I2(1'b0),
    .I3(x39_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011101101001)
) lut_42_30 (
    .O(x42_y30),
    .I0(x40_y27),
    .I1(1'b0),
    .I2(x39_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001100110001)
) lut_43_30 (
    .O(x43_y30),
    .I0(x40_y34),
    .I1(x40_y27),
    .I2(x41_y26),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111100000101)
) lut_44_30 (
    .O(x44_y30),
    .I0(x42_y31),
    .I1(x41_y35),
    .I2(1'b0),
    .I3(x42_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101101110100)
) lut_45_30 (
    .O(x45_y30),
    .I0(x43_y34),
    .I1(x42_y32),
    .I2(1'b0),
    .I3(x42_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011111011111)
) lut_46_30 (
    .O(x46_y30),
    .I0(x44_y27),
    .I1(x44_y35),
    .I2(1'b0),
    .I3(x43_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000101100010)
) lut_47_30 (
    .O(x47_y30),
    .I0(x45_y35),
    .I1(x44_y34),
    .I2(1'b0),
    .I3(x44_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011000110110)
) lut_48_30 (
    .O(x48_y30),
    .I0(x46_y25),
    .I1(x45_y28),
    .I2(x45_y34),
    .I3(x46_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111111101011)
) lut_49_30 (
    .O(x49_y30),
    .I0(1'b0),
    .I1(x47_y27),
    .I2(x46_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111110000101)
) lut_50_30 (
    .O(x50_y30),
    .I0(x48_y25),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x47_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011001001101)
) lut_51_30 (
    .O(x51_y30),
    .I0(x48_y25),
    .I1(1'b0),
    .I2(x48_y28),
    .I3(x48_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111011001000)
) lut_52_30 (
    .O(x52_y30),
    .I0(1'b0),
    .I1(x50_y31),
    .I2(x49_y33),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010100001000)
) lut_53_30 (
    .O(x53_y30),
    .I0(x50_y34),
    .I1(x50_y26),
    .I2(x51_y35),
    .I3(x51_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111011010100)
) lut_54_30 (
    .O(x54_y30),
    .I0(x52_y26),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x52_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110100111100)
) lut_55_30 (
    .O(x55_y30),
    .I0(x53_y35),
    .I1(x52_y27),
    .I2(x52_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101110000000)
) lut_56_30 (
    .O(x56_y30),
    .I0(1'b0),
    .I1(x54_y26),
    .I2(1'b0),
    .I3(x53_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011001011010)
) lut_57_30 (
    .O(x57_y30),
    .I0(x55_y32),
    .I1(x55_y26),
    .I2(x55_y32),
    .I3(x54_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001001001001)
) lut_58_30 (
    .O(x58_y30),
    .I0(1'b0),
    .I1(x55_y29),
    .I2(x56_y29),
    .I3(x55_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100010101011)
) lut_59_30 (
    .O(x59_y30),
    .I0(x57_y35),
    .I1(x56_y34),
    .I2(x56_y28),
    .I3(x56_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000011001010)
) lut_60_30 (
    .O(x60_y30),
    .I0(1'b0),
    .I1(x58_y27),
    .I2(1'b0),
    .I3(x58_y25)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100100100011)
) lut_61_30 (
    .O(x61_y30),
    .I0(1'b0),
    .I1(x58_y29),
    .I2(x58_y25),
    .I3(x58_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011011100011)
) lut_62_30 (
    .O(x62_y30),
    .I0(x59_y33),
    .I1(x60_y33),
    .I2(x60_y32),
    .I3(x60_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000111011001)
) lut_0_31 (
    .O(x0_y31),
    .I0(in1),
    .I1(in3),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001011111101)
) lut_1_31 (
    .O(x1_y31),
    .I0(1'b0),
    .I1(in0),
    .I2(in4),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001111001101)
) lut_2_31 (
    .O(x2_y31),
    .I0(1'b0),
    .I1(in3),
    .I2(in6),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011011110011)
) lut_3_31 (
    .O(x3_y31),
    .I0(in6),
    .I1(x1_y36),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111010001001)
) lut_4_31 (
    .O(x4_y31),
    .I0(x2_y36),
    .I1(x1_y29),
    .I2(x1_y36),
    .I3(x1_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011111011110)
) lut_5_31 (
    .O(x5_y31),
    .I0(x2_y29),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x3_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101101010000)
) lut_6_31 (
    .O(x6_y31),
    .I0(x3_y34),
    .I1(x3_y34),
    .I2(x4_y35),
    .I3(x3_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001111110110)
) lut_7_31 (
    .O(x7_y31),
    .I0(x4_y28),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x5_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000011111100)
) lut_8_31 (
    .O(x8_y31),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x5_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100001000001)
) lut_9_31 (
    .O(x9_y31),
    .I0(x7_y34),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x5_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001001111000)
) lut_10_31 (
    .O(x10_y31),
    .I0(1'b0),
    .I1(x8_y33),
    .I2(x7_y36),
    .I3(x8_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110110001010)
) lut_11_31 (
    .O(x11_y31),
    .I0(x9_y31),
    .I1(x9_y27),
    .I2(x9_y30),
    .I3(x8_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000010001110)
) lut_12_31 (
    .O(x12_y31),
    .I0(x9_y32),
    .I1(x9_y27),
    .I2(x10_y27),
    .I3(x9_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010001001100)
) lut_13_31 (
    .O(x13_y31),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x11_y35),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100001001000)
) lut_14_31 (
    .O(x14_y31),
    .I0(x12_y26),
    .I1(x11_y33),
    .I2(x12_y36),
    .I3(x11_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000111000110)
) lut_15_31 (
    .O(x15_y31),
    .I0(x13_y29),
    .I1(x13_y31),
    .I2(x13_y27),
    .I3(x13_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110110101011)
) lut_16_31 (
    .O(x16_y31),
    .I0(x14_y36),
    .I1(x14_y34),
    .I2(x13_y36),
    .I3(x13_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000101000011)
) lut_17_31 (
    .O(x17_y31),
    .I0(x15_y26),
    .I1(x14_y29),
    .I2(x14_y31),
    .I3(x15_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011011000001)
) lut_18_31 (
    .O(x18_y31),
    .I0(x16_y30),
    .I1(1'b0),
    .I2(x16_y33),
    .I3(x16_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101101100000)
) lut_19_31 (
    .O(x19_y31),
    .I0(x16_y34),
    .I1(1'b0),
    .I2(x17_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010111111011)
) lut_20_31 (
    .O(x20_y31),
    .I0(x18_y27),
    .I1(x17_y34),
    .I2(x18_y27),
    .I3(x17_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110001010010)
) lut_21_31 (
    .O(x21_y31),
    .I0(x18_y35),
    .I1(x18_y36),
    .I2(x18_y28),
    .I3(x19_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001111101000)
) lut_22_31 (
    .O(x22_y31),
    .I0(x20_y33),
    .I1(x20_y35),
    .I2(1'b0),
    .I3(x20_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000001000000)
) lut_23_31 (
    .O(x23_y31),
    .I0(x20_y30),
    .I1(x20_y29),
    .I2(x20_y32),
    .I3(x21_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000011100111)
) lut_24_31 (
    .O(x24_y31),
    .I0(x21_y36),
    .I1(x22_y26),
    .I2(x22_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110011110101)
) lut_25_31 (
    .O(x25_y31),
    .I0(1'b0),
    .I1(x22_y33),
    .I2(1'b0),
    .I3(x22_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010111001101)
) lut_26_31 (
    .O(x26_y31),
    .I0(x23_y29),
    .I1(x23_y33),
    .I2(x23_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110001111101)
) lut_27_31 (
    .O(x27_y31),
    .I0(x24_y35),
    .I1(x24_y30),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001110110100)
) lut_28_31 (
    .O(x28_y31),
    .I0(x26_y27),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x25_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111011011101)
) lut_29_31 (
    .O(x29_y31),
    .I0(x27_y29),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111010110011)
) lut_30_31 (
    .O(x30_y31),
    .I0(1'b0),
    .I1(x27_y36),
    .I2(x27_y26),
    .I3(x27_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011101011010)
) lut_31_31 (
    .O(x31_y31),
    .I0(x28_y33),
    .I1(x29_y28),
    .I2(x28_y33),
    .I3(x28_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011001110101)
) lut_32_31 (
    .O(x32_y31),
    .I0(x29_y27),
    .I1(x30_y30),
    .I2(1'b0),
    .I3(x30_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000000010000)
) lut_33_31 (
    .O(x33_y31),
    .I0(1'b0),
    .I1(x30_y33),
    .I2(x30_y29),
    .I3(x30_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000111000010)
) lut_34_31 (
    .O(x34_y31),
    .I0(x32_y30),
    .I1(x31_y35),
    .I2(x31_y36),
    .I3(x31_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101110000011)
) lut_35_31 (
    .O(x35_y31),
    .I0(x32_y26),
    .I1(x32_y27),
    .I2(1'b0),
    .I3(x32_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100000111111)
) lut_36_31 (
    .O(x36_y31),
    .I0(x33_y34),
    .I1(x33_y36),
    .I2(1'b0),
    .I3(x33_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101111011101)
) lut_37_31 (
    .O(x37_y31),
    .I0(x35_y30),
    .I1(x34_y36),
    .I2(1'b0),
    .I3(x35_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101101111110)
) lut_38_31 (
    .O(x38_y31),
    .I0(x36_y36),
    .I1(x36_y31),
    .I2(x35_y33),
    .I3(x35_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000000110001)
) lut_39_31 (
    .O(x39_y31),
    .I0(x36_y27),
    .I1(x36_y33),
    .I2(x36_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011110101000)
) lut_40_31 (
    .O(x40_y31),
    .I0(x38_y31),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x37_y26)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101001001110)
) lut_41_31 (
    .O(x41_y31),
    .I0(x39_y27),
    .I1(x39_y26),
    .I2(1'b0),
    .I3(x38_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101010100100)
) lut_42_31 (
    .O(x42_y31),
    .I0(x40_y30),
    .I1(1'b0),
    .I2(x40_y36),
    .I3(x39_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100110011000)
) lut_43_31 (
    .O(x43_y31),
    .I0(x40_y28),
    .I1(x40_y33),
    .I2(x40_y33),
    .I3(x40_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111111111011)
) lut_44_31 (
    .O(x44_y31),
    .I0(x41_y28),
    .I1(x41_y26),
    .I2(x42_y29),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100011001001)
) lut_45_31 (
    .O(x45_y31),
    .I0(x42_y31),
    .I1(x43_y31),
    .I2(1'b0),
    .I3(x42_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001000100010)
) lut_46_31 (
    .O(x46_y31),
    .I0(x44_y27),
    .I1(x43_y29),
    .I2(x43_y35),
    .I3(x43_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111011110010)
) lut_47_31 (
    .O(x47_y31),
    .I0(x45_y26),
    .I1(x44_y35),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001101001100)
) lut_48_31 (
    .O(x48_y31),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x46_y27),
    .I3(x45_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001111111100)
) lut_49_31 (
    .O(x49_y31),
    .I0(1'b0),
    .I1(x46_y28),
    .I2(x47_y35),
    .I3(x46_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100110111110)
) lut_50_31 (
    .O(x50_y31),
    .I0(x48_y29),
    .I1(x47_y31),
    .I2(x48_y32),
    .I3(x48_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000111001000)
) lut_51_31 (
    .O(x51_y31),
    .I0(1'b0),
    .I1(x49_y26),
    .I2(x49_y32),
    .I3(x48_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101010001110)
) lut_52_31 (
    .O(x52_y31),
    .I0(x50_y32),
    .I1(x49_y31),
    .I2(x50_y36),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100111010111)
) lut_53_31 (
    .O(x53_y31),
    .I0(1'b0),
    .I1(x51_y26),
    .I2(x50_y31),
    .I3(x51_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101000111001)
) lut_54_31 (
    .O(x54_y31),
    .I0(x51_y26),
    .I1(1'b0),
    .I2(x52_y26),
    .I3(x51_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100000110101)
) lut_55_31 (
    .O(x55_y31),
    .I0(x53_y30),
    .I1(x52_y32),
    .I2(x53_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100101111110)
) lut_56_31 (
    .O(x56_y31),
    .I0(1'b0),
    .I1(x54_y27),
    .I2(x53_y35),
    .I3(x54_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111001101010)
) lut_57_31 (
    .O(x57_y31),
    .I0(x54_y32),
    .I1(x54_y31),
    .I2(x55_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100010000100)
) lut_58_31 (
    .O(x58_y31),
    .I0(x55_y26),
    .I1(x55_y28),
    .I2(x56_y34),
    .I3(x55_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000001101001)
) lut_59_31 (
    .O(x59_y31),
    .I0(x56_y33),
    .I1(x56_y36),
    .I2(1'b0),
    .I3(x57_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010111111010)
) lut_60_31 (
    .O(x60_y31),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x58_y30),
    .I3(x58_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100001000010)
) lut_61_31 (
    .O(x61_y31),
    .I0(x58_y28),
    .I1(x58_y27),
    .I2(x59_y32),
    .I3(x58_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000101100011)
) lut_62_31 (
    .O(x62_y31),
    .I0(x60_y35),
    .I1(x59_y29),
    .I2(1'b0),
    .I3(x60_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011011000011)
) lut_0_32 (
    .O(x0_y32),
    .I0(in2),
    .I1(in2),
    .I2(in6),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001011001010)
) lut_1_32 (
    .O(x1_y32),
    .I0(in2),
    .I1(in3),
    .I2(in8),
    .I3(in9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001011101110)
) lut_2_32 (
    .O(x2_y32),
    .I0(1'b0),
    .I1(in4),
    .I2(in2),
    .I3(in4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010001010110)
) lut_3_32 (
    .O(x3_y32),
    .I0(in4),
    .I1(in4),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010000001011)
) lut_4_32 (
    .O(x4_y32),
    .I0(x2_y35),
    .I1(x1_y29),
    .I2(x1_y27),
    .I3(x2_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001010000001)
) lut_5_32 (
    .O(x5_y32),
    .I0(x3_y32),
    .I1(x2_y37),
    .I2(x2_y36),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000000101110)
) lut_6_32 (
    .O(x6_y32),
    .I0(1'b0),
    .I1(x4_y35),
    .I2(x4_y27),
    .I3(x3_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100101000011)
) lut_7_32 (
    .O(x7_y32),
    .I0(1'b0),
    .I1(x5_y31),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000000111000)
) lut_8_32 (
    .O(x8_y32),
    .I0(x6_y31),
    .I1(x6_y33),
    .I2(x5_y27),
    .I3(x6_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100001101110)
) lut_9_32 (
    .O(x9_y32),
    .I0(x6_y27),
    .I1(1'b0),
    .I2(x5_y27),
    .I3(x6_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100011010110)
) lut_10_32 (
    .O(x10_y32),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x8_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100001111001)
) lut_11_32 (
    .O(x11_y32),
    .I0(x8_y27),
    .I1(1'b0),
    .I2(x9_y32),
    .I3(x8_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010111000000)
) lut_12_32 (
    .O(x12_y32),
    .I0(x10_y28),
    .I1(1'b0),
    .I2(x9_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011010010011)
) lut_13_32 (
    .O(x13_y32),
    .I0(x10_y34),
    .I1(x11_y32),
    .I2(1'b0),
    .I3(x11_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000000011100)
) lut_14_32 (
    .O(x14_y32),
    .I0(x12_y37),
    .I1(x12_y35),
    .I2(x11_y34),
    .I3(x12_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110011011011)
) lut_15_32 (
    .O(x15_y32),
    .I0(x12_y29),
    .I1(x13_y27),
    .I2(x12_y36),
    .I3(x12_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000001100100)
) lut_16_32 (
    .O(x16_y32),
    .I0(x14_y28),
    .I1(1'b0),
    .I2(x14_y27),
    .I3(x14_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010110101110)
) lut_17_32 (
    .O(x17_y32),
    .I0(x14_y37),
    .I1(x15_y27),
    .I2(1'b0),
    .I3(x15_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101100100010)
) lut_18_32 (
    .O(x18_y32),
    .I0(x15_y36),
    .I1(1'b0),
    .I2(x15_y29),
    .I3(x15_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011000000001)
) lut_19_32 (
    .O(x19_y32),
    .I0(x16_y29),
    .I1(1'b0),
    .I2(x17_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010101001010)
) lut_20_32 (
    .O(x20_y32),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101111100100)
) lut_21_32 (
    .O(x21_y32),
    .I0(x18_y37),
    .I1(1'b0),
    .I2(x19_y37),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110101111110)
) lut_22_32 (
    .O(x22_y32),
    .I0(x19_y29),
    .I1(x20_y27),
    .I2(x19_y30),
    .I3(x19_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101111101000)
) lut_23_32 (
    .O(x23_y32),
    .I0(1'b0),
    .I1(x20_y29),
    .I2(x21_y35),
    .I3(x21_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110100010011)
) lut_24_32 (
    .O(x24_y32),
    .I0(x21_y28),
    .I1(x21_y27),
    .I2(1'b0),
    .I3(x22_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001111110100)
) lut_25_32 (
    .O(x25_y32),
    .I0(x23_y36),
    .I1(x22_y33),
    .I2(x23_y33),
    .I3(x22_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110010010101)
) lut_26_32 (
    .O(x26_y32),
    .I0(x24_y35),
    .I1(x23_y30),
    .I2(x23_y27),
    .I3(x23_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101010110110)
) lut_27_32 (
    .O(x27_y32),
    .I0(1'b0),
    .I1(x25_y27),
    .I2(x24_y35),
    .I3(x24_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110001011001)
) lut_28_32 (
    .O(x28_y32),
    .I0(x26_y35),
    .I1(x25_y35),
    .I2(x25_y29),
    .I3(x26_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101101110100)
) lut_29_32 (
    .O(x29_y32),
    .I0(x27_y32),
    .I1(1'b0),
    .I2(x27_y29),
    .I3(x26_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011010100100)
) lut_30_32 (
    .O(x30_y32),
    .I0(x28_y34),
    .I1(x28_y37),
    .I2(x27_y36),
    .I3(x27_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010101010010)
) lut_31_32 (
    .O(x31_y32),
    .I0(1'b0),
    .I1(x29_y27),
    .I2(x28_y31),
    .I3(x29_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110110011011)
) lut_32_32 (
    .O(x32_y32),
    .I0(x29_y29),
    .I1(x29_y37),
    .I2(x30_y30),
    .I3(x29_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010100011011)
) lut_33_32 (
    .O(x33_y32),
    .I0(1'b0),
    .I1(x31_y29),
    .I2(x31_y33),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100101100111)
) lut_34_32 (
    .O(x34_y32),
    .I0(x31_y33),
    .I1(1'b0),
    .I2(x32_y28),
    .I3(x32_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000100101110)
) lut_35_32 (
    .O(x35_y32),
    .I0(x33_y36),
    .I1(x32_y32),
    .I2(x32_y35),
    .I3(x32_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011100100111)
) lut_36_32 (
    .O(x36_y32),
    .I0(1'b0),
    .I1(x33_y37),
    .I2(x34_y34),
    .I3(x34_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110101010101)
) lut_37_32 (
    .O(x37_y32),
    .I0(x34_y33),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x35_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000111110101)
) lut_38_32 (
    .O(x38_y32),
    .I0(1'b0),
    .I1(x36_y32),
    .I2(1'b0),
    .I3(x35_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010010001001)
) lut_39_32 (
    .O(x39_y32),
    .I0(1'b0),
    .I1(x37_y27),
    .I2(x37_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000000100011)
) lut_40_32 (
    .O(x40_y32),
    .I0(x37_y35),
    .I1(1'b0),
    .I2(x38_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111101000000)
) lut_41_32 (
    .O(x41_y32),
    .I0(1'b0),
    .I1(x39_y29),
    .I2(x39_y37),
    .I3(x39_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110011011101)
) lut_42_32 (
    .O(x42_y32),
    .I0(x40_y33),
    .I1(x39_y35),
    .I2(x39_y29),
    .I3(x39_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000010011110)
) lut_43_32 (
    .O(x43_y32),
    .I0(x41_y31),
    .I1(x41_y36),
    .I2(x40_y33),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100010011110)
) lut_44_32 (
    .O(x44_y32),
    .I0(1'b0),
    .I1(x42_y34),
    .I2(1'b0),
    .I3(x42_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000110011000)
) lut_45_32 (
    .O(x45_y32),
    .I0(1'b0),
    .I1(x42_y34),
    .I2(x42_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000100110100)
) lut_46_32 (
    .O(x46_y32),
    .I0(x44_y32),
    .I1(x44_y31),
    .I2(x43_y30),
    .I3(x43_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000000110011)
) lut_47_32 (
    .O(x47_y32),
    .I0(x45_y37),
    .I1(x44_y30),
    .I2(1'b0),
    .I3(x45_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111001010010)
) lut_48_32 (
    .O(x48_y32),
    .I0(x46_y31),
    .I1(x46_y30),
    .I2(x46_y35),
    .I3(x46_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011111001111)
) lut_49_32 (
    .O(x49_y32),
    .I0(x46_y36),
    .I1(x47_y28),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111000001100)
) lut_50_32 (
    .O(x50_y32),
    .I0(x48_y29),
    .I1(x47_y33),
    .I2(x47_y34),
    .I3(x47_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010011111010)
) lut_51_32 (
    .O(x51_y32),
    .I0(1'b0),
    .I1(x49_y29),
    .I2(x48_y30),
    .I3(x48_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111010011101)
) lut_52_32 (
    .O(x52_y32),
    .I0(x50_y33),
    .I1(1'b0),
    .I2(x49_y30),
    .I3(x50_y27)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010101110011)
) lut_53_32 (
    .O(x53_y32),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x50_y37),
    .I3(x50_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101111110101)
) lut_54_32 (
    .O(x54_y32),
    .I0(1'b0),
    .I1(x52_y31),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110001110000)
) lut_55_32 (
    .O(x55_y32),
    .I0(x52_y28),
    .I1(1'b0),
    .I2(x53_y31),
    .I3(x52_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101001000001)
) lut_56_32 (
    .O(x56_y32),
    .I0(x54_y30),
    .I1(x54_y36),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011101110011)
) lut_57_32 (
    .O(x57_y32),
    .I0(x55_y29),
    .I1(x54_y37),
    .I2(x55_y35),
    .I3(x54_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101101011100)
) lut_58_32 (
    .O(x58_y32),
    .I0(x55_y29),
    .I1(x56_y28),
    .I2(x56_y34),
    .I3(x55_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011110110010)
) lut_59_32 (
    .O(x59_y32),
    .I0(x56_y32),
    .I1(x57_y32),
    .I2(x56_y35),
    .I3(x57_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111111010010)
) lut_60_32 (
    .O(x60_y32),
    .I0(x58_y27),
    .I1(x57_y33),
    .I2(x57_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101111110110)
) lut_61_32 (
    .O(x61_y32),
    .I0(x59_y32),
    .I1(x59_y30),
    .I2(x58_y33),
    .I3(x58_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001111110100)
) lut_62_32 (
    .O(x62_y32),
    .I0(1'b0),
    .I1(x60_y34),
    .I2(x60_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000110001111)
) lut_0_33 (
    .O(x0_y33),
    .I0(in7),
    .I1(in8),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100000000100)
) lut_1_33 (
    .O(x1_y33),
    .I0(in4),
    .I1(in9),
    .I2(in7),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011011011000)
) lut_2_33 (
    .O(x2_y33),
    .I0(in7),
    .I1(in8),
    .I2(in0),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111011101100)
) lut_3_33 (
    .O(x3_y33),
    .I0(x1_y33),
    .I1(1'b0),
    .I2(in5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101111101110)
) lut_4_33 (
    .O(x4_y33),
    .I0(1'b0),
    .I1(x2_y28),
    .I2(x2_y31),
    .I3(x1_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010010100110)
) lut_5_33 (
    .O(x5_y33),
    .I0(x2_y31),
    .I1(x2_y29),
    .I2(1'b0),
    .I3(x3_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100010010110)
) lut_6_33 (
    .O(x6_y33),
    .I0(1'b0),
    .I1(x4_y29),
    .I2(x3_y35),
    .I3(x4_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001000101101)
) lut_7_33 (
    .O(x7_y33),
    .I0(1'b0),
    .I1(x4_y38),
    .I2(x5_y37),
    .I3(x4_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010010000000)
) lut_8_33 (
    .O(x8_y33),
    .I0(1'b0),
    .I1(x6_y33),
    .I2(x5_y31),
    .I3(x6_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011110101111)
) lut_9_33 (
    .O(x9_y33),
    .I0(x6_y38),
    .I1(1'b0),
    .I2(x5_y31),
    .I3(x6_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010110000000)
) lut_10_33 (
    .O(x10_y33),
    .I0(x8_y31),
    .I1(x7_y33),
    .I2(1'b0),
    .I3(x8_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000001010100)
) lut_11_33 (
    .O(x11_y33),
    .I0(x8_y35),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x8_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001101011110)
) lut_12_33 (
    .O(x12_y33),
    .I0(x9_y38),
    .I1(x9_y38),
    .I2(x10_y35),
    .I3(x10_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001010011001)
) lut_13_33 (
    .O(x13_y33),
    .I0(x11_y38),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x11_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100100111000)
) lut_14_33 (
    .O(x14_y33),
    .I0(x12_y34),
    .I1(1'b0),
    .I2(x11_y29),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100100000011)
) lut_15_33 (
    .O(x15_y33),
    .I0(x12_y28),
    .I1(1'b0),
    .I2(x12_y36),
    .I3(x13_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110110101001)
) lut_16_33 (
    .O(x16_y33),
    .I0(x13_y35),
    .I1(x13_y33),
    .I2(x13_y35),
    .I3(x14_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110000011001)
) lut_17_33 (
    .O(x17_y33),
    .I0(x15_y28),
    .I1(x14_y32),
    .I2(1'b0),
    .I3(x14_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110010101110)
) lut_18_33 (
    .O(x18_y33),
    .I0(1'b0),
    .I1(x16_y28),
    .I2(x16_y35),
    .I3(x16_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010010001001)
) lut_19_33 (
    .O(x19_y33),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x16_y32),
    .I3(x17_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110101100010)
) lut_20_33 (
    .O(x20_y33),
    .I0(x18_y32),
    .I1(x17_y32),
    .I2(x17_y31),
    .I3(x17_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110110101110)
) lut_21_33 (
    .O(x21_y33),
    .I0(1'b0),
    .I1(x18_y33),
    .I2(1'b0),
    .I3(x18_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110110010111)
) lut_22_33 (
    .O(x22_y33),
    .I0(x19_y30),
    .I1(x19_y28),
    .I2(x20_y38),
    .I3(x19_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111011100111)
) lut_23_33 (
    .O(x23_y33),
    .I0(1'b0),
    .I1(x21_y37),
    .I2(x21_y31),
    .I3(x20_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110000110100)
) lut_24_33 (
    .O(x24_y33),
    .I0(x21_y31),
    .I1(x21_y35),
    .I2(x22_y31),
    .I3(x22_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111110100001)
) lut_25_33 (
    .O(x25_y33),
    .I0(x22_y29),
    .I1(x22_y30),
    .I2(x22_y35),
    .I3(x23_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110001100101)
) lut_26_33 (
    .O(x26_y33),
    .I0(x23_y34),
    .I1(1'b0),
    .I2(x23_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101110110110)
) lut_27_33 (
    .O(x27_y33),
    .I0(x25_y35),
    .I1(x24_y35),
    .I2(x24_y34),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011000101011)
) lut_28_33 (
    .O(x28_y33),
    .I0(x26_y32),
    .I1(x25_y32),
    .I2(x26_y37),
    .I3(x25_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100110110110)
) lut_29_33 (
    .O(x29_y33),
    .I0(x27_y36),
    .I1(x27_y32),
    .I2(1'b0),
    .I3(x27_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100001101000)
) lut_30_33 (
    .O(x30_y33),
    .I0(x28_y28),
    .I1(x28_y31),
    .I2(x28_y38),
    .I3(x27_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100001011110)
) lut_31_33 (
    .O(x31_y33),
    .I0(1'b0),
    .I1(x29_y29),
    .I2(x29_y36),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010110110011)
) lut_32_33 (
    .O(x32_y33),
    .I0(1'b0),
    .I1(x29_y36),
    .I2(x29_y30),
    .I3(x29_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001110110001)
) lut_33_33 (
    .O(x33_y33),
    .I0(x31_y28),
    .I1(1'b0),
    .I2(x30_y28),
    .I3(x31_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100101001011)
) lut_34_33 (
    .O(x34_y33),
    .I0(1'b0),
    .I1(x31_y36),
    .I2(1'b0),
    .I3(x31_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101010000111)
) lut_35_33 (
    .O(x35_y33),
    .I0(x32_y28),
    .I1(1'b0),
    .I2(x32_y36),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000001001011)
) lut_36_33 (
    .O(x36_y33),
    .I0(x34_y29),
    .I1(x33_y36),
    .I2(x34_y31),
    .I3(x33_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010001000001)
) lut_37_33 (
    .O(x37_y33),
    .I0(1'b0),
    .I1(x35_y34),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100100011011)
) lut_38_33 (
    .O(x38_y33),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x35_y36),
    .I3(x35_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101100101011)
) lut_39_33 (
    .O(x39_y33),
    .I0(x37_y37),
    .I1(x37_y31),
    .I2(x37_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000100001000)
) lut_40_33 (
    .O(x40_y33),
    .I0(1'b0),
    .I1(x38_y28),
    .I2(x37_y37),
    .I3(x38_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010000000010)
) lut_41_33 (
    .O(x41_y33),
    .I0(x39_y28),
    .I1(x38_y32),
    .I2(x38_y38),
    .I3(x38_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001000010111)
) lut_42_33 (
    .O(x42_y33),
    .I0(x40_y30),
    .I1(x40_y31),
    .I2(x39_y35),
    .I3(x39_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001011110110)
) lut_43_33 (
    .O(x43_y33),
    .I0(1'b0),
    .I1(x41_y33),
    .I2(x41_y28),
    .I3(x40_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011110110000)
) lut_44_33 (
    .O(x44_y33),
    .I0(x41_y34),
    .I1(x42_y30),
    .I2(x42_y38),
    .I3(x42_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010101100101)
) lut_45_33 (
    .O(x45_y33),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x43_y30),
    .I3(x43_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111001111100)
) lut_46_33 (
    .O(x46_y33),
    .I0(x44_y35),
    .I1(x43_y31),
    .I2(x44_y30),
    .I3(x43_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110101011001)
) lut_47_33 (
    .O(x47_y33),
    .I0(x45_y32),
    .I1(x45_y37),
    .I2(x44_y32),
    .I3(x44_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010010011011)
) lut_48_33 (
    .O(x48_y33),
    .I0(x46_y29),
    .I1(x45_y38),
    .I2(x45_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110001001010)
) lut_49_33 (
    .O(x49_y33),
    .I0(x46_y34),
    .I1(x47_y34),
    .I2(x46_y29),
    .I3(x46_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100011101110)
) lut_50_33 (
    .O(x50_y33),
    .I0(x47_y29),
    .I1(1'b0),
    .I2(x47_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000001010000)
) lut_51_33 (
    .O(x51_y33),
    .I0(x49_y35),
    .I1(x49_y33),
    .I2(x49_y36),
    .I3(x49_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011100111000)
) lut_52_33 (
    .O(x52_y33),
    .I0(x49_y34),
    .I1(x49_y34),
    .I2(1'b0),
    .I3(x50_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010111000110)
) lut_53_33 (
    .O(x53_y33),
    .I0(x50_y37),
    .I1(x50_y33),
    .I2(x51_y37),
    .I3(x51_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010110010101)
) lut_54_33 (
    .O(x54_y33),
    .I0(x51_y38),
    .I1(x52_y38),
    .I2(x51_y34),
    .I3(x52_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010001110010)
) lut_55_33 (
    .O(x55_y33),
    .I0(x52_y31),
    .I1(x53_y30),
    .I2(1'b0),
    .I3(x52_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110111010110)
) lut_56_33 (
    .O(x56_y33),
    .I0(x53_y31),
    .I1(x54_y30),
    .I2(x53_y31),
    .I3(x54_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001111000100)
) lut_57_33 (
    .O(x57_y33),
    .I0(x54_y32),
    .I1(x55_y37),
    .I2(x55_y36),
    .I3(x54_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101101000110)
) lut_58_33 (
    .O(x58_y33),
    .I0(x56_y30),
    .I1(1'b0),
    .I2(x55_y32),
    .I3(x56_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000101011011)
) lut_59_33 (
    .O(x59_y33),
    .I0(x57_y30),
    .I1(x57_y36),
    .I2(x57_y28),
    .I3(x56_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001111101010)
) lut_60_33 (
    .O(x60_y33),
    .I0(x58_y37),
    .I1(1'b0),
    .I2(x57_y38),
    .I3(x57_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111011010101)
) lut_61_33 (
    .O(x61_y33),
    .I0(x58_y37),
    .I1(x59_y31),
    .I2(x58_y37),
    .I3(x59_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001010101011)
) lut_62_33 (
    .O(x62_y33),
    .I0(x60_y31),
    .I1(x60_y30),
    .I2(x60_y35),
    .I3(x60_y28)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000100101010)
) lut_0_34 (
    .O(x0_y34),
    .I0(in3),
    .I1(in6),
    .I2(in9),
    .I3(in1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100100110111)
) lut_1_34 (
    .O(x1_y34),
    .I0(in4),
    .I1(in7),
    .I2(in2),
    .I3(in9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100000010011)
) lut_2_34 (
    .O(x2_y34),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111101111010)
) lut_3_34 (
    .O(x3_y34),
    .I0(in5),
    .I1(1'b0),
    .I2(x1_y35),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010100111100)
) lut_4_34 (
    .O(x4_y34),
    .I0(x2_y38),
    .I1(x2_y34),
    .I2(x2_y39),
    .I3(x2_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101000011110)
) lut_5_34 (
    .O(x5_y34),
    .I0(x2_y33),
    .I1(x3_y31),
    .I2(x2_y36),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111010110010)
) lut_6_34 (
    .O(x6_y34),
    .I0(x4_y35),
    .I1(x4_y36),
    .I2(x4_y38),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011011111100)
) lut_7_34 (
    .O(x7_y34),
    .I0(x4_y38),
    .I1(1'b0),
    .I2(x4_y32),
    .I3(x5_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111011001000)
) lut_8_34 (
    .O(x8_y34),
    .I0(1'b0),
    .I1(x5_y34),
    .I2(x6_y30),
    .I3(x5_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000110001010)
) lut_9_34 (
    .O(x9_y34),
    .I0(x6_y36),
    .I1(x7_y30),
    .I2(x6_y30),
    .I3(x5_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100100101001)
) lut_10_34 (
    .O(x10_y34),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x7_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110000110000)
) lut_11_34 (
    .O(x11_y34),
    .I0(x9_y33),
    .I1(x8_y30),
    .I2(1'b0),
    .I3(x9_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001010100010)
) lut_12_34 (
    .O(x12_y34),
    .I0(x10_y30),
    .I1(x10_y30),
    .I2(x10_y35),
    .I3(x9_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010001000101)
) lut_13_34 (
    .O(x13_y34),
    .I0(x11_y39),
    .I1(x11_y30),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100110001110)
) lut_14_34 (
    .O(x14_y34),
    .I0(x11_y33),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x11_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011011001101)
) lut_15_34 (
    .O(x15_y34),
    .I0(x13_y29),
    .I1(x12_y31),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001110001001)
) lut_16_34 (
    .O(x16_y34),
    .I0(x13_y36),
    .I1(x13_y29),
    .I2(x13_y39),
    .I3(x14_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100010001000)
) lut_17_34 (
    .O(x17_y34),
    .I0(1'b0),
    .I1(x15_y36),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000011011110)
) lut_18_34 (
    .O(x18_y34),
    .I0(x15_y39),
    .I1(1'b0),
    .I2(x16_y34),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011011010111)
) lut_19_34 (
    .O(x19_y34),
    .I0(x16_y33),
    .I1(x16_y36),
    .I2(x17_y33),
    .I3(x17_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111010111110)
) lut_20_34 (
    .O(x20_y34),
    .I0(1'b0),
    .I1(x17_y38),
    .I2(1'b0),
    .I3(x17_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001101000011)
) lut_21_34 (
    .O(x21_y34),
    .I0(1'b0),
    .I1(x19_y30),
    .I2(x19_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110110010000)
) lut_22_34 (
    .O(x22_y34),
    .I0(x19_y31),
    .I1(1'b0),
    .I2(x20_y30),
    .I3(x20_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100110110100)
) lut_23_34 (
    .O(x23_y34),
    .I0(x21_y33),
    .I1(x20_y31),
    .I2(x21_y36),
    .I3(x20_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100000110100)
) lut_24_34 (
    .O(x24_y34),
    .I0(1'b0),
    .I1(x21_y35),
    .I2(x21_y30),
    .I3(x21_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100011001011)
) lut_25_34 (
    .O(x25_y34),
    .I0(1'b0),
    .I1(x23_y32),
    .I2(x22_y38),
    .I3(x22_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001011000010)
) lut_26_34 (
    .O(x26_y34),
    .I0(x23_y36),
    .I1(1'b0),
    .I2(x24_y33),
    .I3(x24_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001101100011)
) lut_27_34 (
    .O(x27_y34),
    .I0(1'b0),
    .I1(x24_y35),
    .I2(x25_y33),
    .I3(x25_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101011000011)
) lut_28_34 (
    .O(x28_y34),
    .I0(1'b0),
    .I1(x25_y30),
    .I2(x25_y32),
    .I3(x26_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111011000111)
) lut_29_34 (
    .O(x29_y34),
    .I0(x27_y30),
    .I1(x27_y38),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001000011111)
) lut_30_34 (
    .O(x30_y34),
    .I0(1'b0),
    .I1(x28_y29),
    .I2(x27_y32),
    .I3(x27_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101100111110)
) lut_31_34 (
    .O(x31_y34),
    .I0(x28_y39),
    .I1(x28_y36),
    .I2(x28_y32),
    .I3(x28_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011100011001)
) lut_32_34 (
    .O(x32_y34),
    .I0(1'b0),
    .I1(x30_y39),
    .I2(x29_y32),
    .I3(x30_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010010110011)
) lut_33_34 (
    .O(x33_y34),
    .I0(x30_y36),
    .I1(x31_y29),
    .I2(x31_y29),
    .I3(x30_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111101101110)
) lut_34_34 (
    .O(x34_y34),
    .I0(x32_y31),
    .I1(x31_y35),
    .I2(1'b0),
    .I3(x31_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101100111001)
) lut_35_34 (
    .O(x35_y34),
    .I0(x32_y39),
    .I1(x32_y32),
    .I2(x32_y38),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100100000010)
) lut_36_34 (
    .O(x36_y34),
    .I0(x33_y38),
    .I1(x33_y36),
    .I2(1'b0),
    .I3(x34_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111111101110)
) lut_37_34 (
    .O(x37_y34),
    .I0(x34_y33),
    .I1(x34_y34),
    .I2(x34_y36),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011110011111)
) lut_38_34 (
    .O(x38_y34),
    .I0(x36_y31),
    .I1(x35_y33),
    .I2(x35_y38),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100010001101)
) lut_39_34 (
    .O(x39_y34),
    .I0(x36_y39),
    .I1(x37_y32),
    .I2(x37_y30),
    .I3(x37_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010100101010)
) lut_40_34 (
    .O(x40_y34),
    .I0(x37_y33),
    .I1(x37_y35),
    .I2(x38_y32),
    .I3(x38_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001110111011)
) lut_41_34 (
    .O(x41_y34),
    .I0(1'b0),
    .I1(x38_y29),
    .I2(x38_y36),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101110101111)
) lut_42_34 (
    .O(x42_y34),
    .I0(x39_y31),
    .I1(x39_y29),
    .I2(x40_y34),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000101111110)
) lut_43_34 (
    .O(x43_y34),
    .I0(x41_y32),
    .I1(x40_y37),
    .I2(x41_y34),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101100010000)
) lut_44_34 (
    .O(x44_y34),
    .I0(x42_y29),
    .I1(1'b0),
    .I2(x42_y29),
    .I3(x41_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010100101010)
) lut_45_34 (
    .O(x45_y34),
    .I0(x42_y30),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101011101010)
) lut_46_34 (
    .O(x46_y34),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x44_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010110110100)
) lut_47_34 (
    .O(x47_y34),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x44_y32),
    .I3(x45_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111001000011)
) lut_48_34 (
    .O(x48_y34),
    .I0(x45_y32),
    .I1(x46_y29),
    .I2(x46_y35),
    .I3(x45_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100011100011)
) lut_49_34 (
    .O(x49_y34),
    .I0(x46_y35),
    .I1(x46_y33),
    .I2(x46_y35),
    .I3(x47_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110011110110)
) lut_50_34 (
    .O(x50_y34),
    .I0(1'b0),
    .I1(x48_y38),
    .I2(1'b0),
    .I3(x47_y29)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011001011001)
) lut_51_34 (
    .O(x51_y34),
    .I0(x48_y38),
    .I1(x49_y31),
    .I2(x49_y29),
    .I3(x49_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011110001110)
) lut_52_34 (
    .O(x52_y34),
    .I0(x50_y30),
    .I1(x50_y38),
    .I2(x49_y31),
    .I3(x50_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001101110101)
) lut_53_34 (
    .O(x53_y34),
    .I0(x50_y31),
    .I1(x50_y31),
    .I2(x51_y37),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000010010011)
) lut_54_34 (
    .O(x54_y34),
    .I0(1'b0),
    .I1(x52_y38),
    .I2(x52_y29),
    .I3(x52_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000101010010)
) lut_55_34 (
    .O(x55_y34),
    .I0(1'b0),
    .I1(x52_y35),
    .I2(x52_y38),
    .I3(x53_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101011100001)
) lut_56_34 (
    .O(x56_y34),
    .I0(x54_y35),
    .I1(x53_y35),
    .I2(x54_y30),
    .I3(x54_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101110001000)
) lut_57_34 (
    .O(x57_y34),
    .I0(1'b0),
    .I1(x54_y39),
    .I2(x55_y31),
    .I3(x55_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111100000001)
) lut_58_34 (
    .O(x58_y34),
    .I0(x56_y34),
    .I1(x56_y32),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101001100011)
) lut_59_34 (
    .O(x59_y34),
    .I0(x56_y30),
    .I1(x57_y35),
    .I2(x56_y29),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011101101110)
) lut_60_34 (
    .O(x60_y34),
    .I0(x58_y37),
    .I1(x58_y36),
    .I2(x57_y33),
    .I3(x57_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111111111010)
) lut_61_34 (
    .O(x61_y34),
    .I0(x58_y30),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101001101100)
) lut_62_34 (
    .O(x62_y34),
    .I0(x59_y39),
    .I1(1'b0),
    .I2(x60_y39),
    .I3(x59_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100000011010)
) lut_0_35 (
    .O(x0_y35),
    .I0(in8),
    .I1(in0),
    .I2(in3),
    .I3(in9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111110010001)
) lut_1_35 (
    .O(x1_y35),
    .I0(in4),
    .I1(in9),
    .I2(1'b0),
    .I3(in4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010110111000)
) lut_2_35 (
    .O(x2_y35),
    .I0(1'b0),
    .I1(in5),
    .I2(in6),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011100000100)
) lut_3_35 (
    .O(x3_y35),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x1_y33),
    .I3(x1_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000010110111)
) lut_4_35 (
    .O(x4_y35),
    .I0(1'b0),
    .I1(x2_y36),
    .I2(x2_y33),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100011011011)
) lut_5_35 (
    .O(x5_y35),
    .I0(x2_y34),
    .I1(x2_y35),
    .I2(1'b0),
    .I3(x2_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000100001011)
) lut_6_35 (
    .O(x6_y35),
    .I0(x3_y37),
    .I1(x4_y36),
    .I2(x3_y35),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111011011011)
) lut_7_35 (
    .O(x7_y35),
    .I0(x4_y33),
    .I1(x5_y33),
    .I2(x5_y35),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101111011101)
) lut_8_35 (
    .O(x8_y35),
    .I0(x5_y37),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x6_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011010010100)
) lut_9_35 (
    .O(x9_y35),
    .I0(x7_y38),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x6_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111010010011)
) lut_10_35 (
    .O(x10_y35),
    .I0(x8_y38),
    .I1(x7_y35),
    .I2(x8_y38),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001111110100)
) lut_11_35 (
    .O(x11_y35),
    .I0(1'b0),
    .I1(x9_y35),
    .I2(x8_y38),
    .I3(x8_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001010001111)
) lut_12_35 (
    .O(x12_y35),
    .I0(x9_y30),
    .I1(x10_y35),
    .I2(x10_y37),
    .I3(x10_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110101010100)
) lut_13_35 (
    .O(x13_y35),
    .I0(x11_y37),
    .I1(x11_y34),
    .I2(1'b0),
    .I3(x10_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011010100110)
) lut_14_35 (
    .O(x14_y35),
    .I0(x11_y31),
    .I1(x11_y39),
    .I2(x12_y37),
    .I3(x11_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111001001111)
) lut_15_35 (
    .O(x15_y35),
    .I0(x12_y34),
    .I1(x12_y38),
    .I2(x13_y30),
    .I3(x12_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100101101000)
) lut_16_35 (
    .O(x16_y35),
    .I0(1'b0),
    .I1(x14_y34),
    .I2(1'b0),
    .I3(x13_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100010011101)
) lut_17_35 (
    .O(x17_y35),
    .I0(x14_y40),
    .I1(x15_y39),
    .I2(1'b0),
    .I3(x14_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000011110011)
) lut_18_35 (
    .O(x18_y35),
    .I0(1'b0),
    .I1(x15_y34),
    .I2(x15_y33),
    .I3(x15_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111100010011)
) lut_19_35 (
    .O(x19_y35),
    .I0(x17_y33),
    .I1(x16_y31),
    .I2(x16_y33),
    .I3(x16_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011011010101)
) lut_20_35 (
    .O(x20_y35),
    .I0(x17_y38),
    .I1(1'b0),
    .I2(x18_y35),
    .I3(x17_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011000001011)
) lut_21_35 (
    .O(x21_y35),
    .I0(x18_y39),
    .I1(x18_y39),
    .I2(x18_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100111000010)
) lut_22_35 (
    .O(x22_y35),
    .I0(x19_y35),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x19_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000101011000)
) lut_23_35 (
    .O(x23_y35),
    .I0(1'b0),
    .I1(x20_y31),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110111101000)
) lut_24_35 (
    .O(x24_y35),
    .I0(x22_y33),
    .I1(1'b0),
    .I2(x22_y30),
    .I3(x22_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110010110101)
) lut_25_35 (
    .O(x25_y35),
    .I0(x23_y40),
    .I1(x22_y40),
    .I2(x22_y36),
    .I3(x22_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111111011011)
) lut_26_35 (
    .O(x26_y35),
    .I0(1'b0),
    .I1(x23_y30),
    .I2(x24_y33),
    .I3(x23_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100101110000)
) lut_27_35 (
    .O(x27_y35),
    .I0(x24_y37),
    .I1(x25_y37),
    .I2(x25_y33),
    .I3(x24_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000111100001)
) lut_28_35 (
    .O(x28_y35),
    .I0(x26_y36),
    .I1(x25_y34),
    .I2(x26_y37),
    .I3(x26_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111010110011)
) lut_29_35 (
    .O(x29_y35),
    .I0(x26_y39),
    .I1(x27_y34),
    .I2(x26_y39),
    .I3(x27_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000101111011)
) lut_30_35 (
    .O(x30_y35),
    .I0(x28_y39),
    .I1(x28_y35),
    .I2(x28_y39),
    .I3(x27_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111100000100)
) lut_31_35 (
    .O(x31_y35),
    .I0(x29_y38),
    .I1(x28_y31),
    .I2(x28_y39),
    .I3(x29_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010010101110)
) lut_32_35 (
    .O(x32_y35),
    .I0(x29_y38),
    .I1(1'b0),
    .I2(x30_y35),
    .I3(x29_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000001110001)
) lut_33_35 (
    .O(x33_y35),
    .I0(x30_y38),
    .I1(1'b0),
    .I2(x31_y35),
    .I3(x30_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001001101010)
) lut_34_35 (
    .O(x34_y35),
    .I0(x32_y32),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x31_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001001100000)
) lut_35_35 (
    .O(x35_y35),
    .I0(1'b0),
    .I1(x33_y36),
    .I2(x33_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101100111010)
) lut_36_35 (
    .O(x36_y35),
    .I0(x33_y37),
    .I1(x33_y38),
    .I2(x33_y38),
    .I3(x33_y30)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011010110011)
) lut_37_35 (
    .O(x37_y35),
    .I0(x34_y40),
    .I1(x34_y39),
    .I2(x35_y30),
    .I3(x34_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111010011100)
) lut_38_35 (
    .O(x38_y35),
    .I0(x35_y38),
    .I1(1'b0),
    .I2(x36_y33),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101100101011)
) lut_39_35 (
    .O(x39_y35),
    .I0(x36_y36),
    .I1(x37_y40),
    .I2(x37_y37),
    .I3(x36_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010001011001)
) lut_40_35 (
    .O(x40_y35),
    .I0(x38_y38),
    .I1(x38_y35),
    .I2(x37_y33),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000111100111)
) lut_41_35 (
    .O(x41_y35),
    .I0(x38_y30),
    .I1(1'b0),
    .I2(x38_y34),
    .I3(x39_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010100000100)
) lut_42_35 (
    .O(x42_y35),
    .I0(x40_y36),
    .I1(x39_y33),
    .I2(x40_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101110000000)
) lut_43_35 (
    .O(x43_y35),
    .I0(x41_y34),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x41_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110110000000)
) lut_44_35 (
    .O(x44_y35),
    .I0(x41_y34),
    .I1(x41_y31),
    .I2(1'b0),
    .I3(x42_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011001110100)
) lut_45_35 (
    .O(x45_y35),
    .I0(x43_y33),
    .I1(1'b0),
    .I2(x42_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000011110001)
) lut_46_35 (
    .O(x46_y35),
    .I0(x44_y36),
    .I1(x43_y34),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111011100110)
) lut_47_35 (
    .O(x47_y35),
    .I0(x45_y31),
    .I1(x45_y40),
    .I2(x45_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010100001110)
) lut_48_35 (
    .O(x48_y35),
    .I0(1'b0),
    .I1(x46_y40),
    .I2(x46_y32),
    .I3(x45_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010111111001)
) lut_49_35 (
    .O(x49_y35),
    .I0(x46_y37),
    .I1(x47_y38),
    .I2(x47_y33),
    .I3(x46_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111100100111)
) lut_50_35 (
    .O(x50_y35),
    .I0(x48_y34),
    .I1(x48_y36),
    .I2(x48_y32),
    .I3(x48_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001000111110)
) lut_51_35 (
    .O(x51_y35),
    .I0(x48_y39),
    .I1(x49_y32),
    .I2(x48_y38),
    .I3(x49_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111110111011)
) lut_52_35 (
    .O(x52_y35),
    .I0(1'b0),
    .I1(x50_y36),
    .I2(1'b0),
    .I3(x50_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001010111001)
) lut_53_35 (
    .O(x53_y35),
    .I0(x51_y35),
    .I1(x51_y39),
    .I2(x50_y37),
    .I3(x50_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110010110011)
) lut_54_35 (
    .O(x54_y35),
    .I0(x51_y37),
    .I1(x51_y31),
    .I2(x51_y35),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111000000111)
) lut_55_35 (
    .O(x55_y35),
    .I0(x53_y38),
    .I1(x52_y31),
    .I2(x52_y30),
    .I3(x52_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000010111100)
) lut_56_35 (
    .O(x56_y35),
    .I0(x54_y34),
    .I1(x53_y34),
    .I2(x53_y37),
    .I3(x54_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011000011000)
) lut_57_35 (
    .O(x57_y35),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x54_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000010001111)
) lut_58_35 (
    .O(x58_y35),
    .I0(x55_y32),
    .I1(x55_y35),
    .I2(x55_y34),
    .I3(x55_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101100111001)
) lut_59_35 (
    .O(x59_y35),
    .I0(x57_y38),
    .I1(x57_y37),
    .I2(x56_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000000101111)
) lut_60_35 (
    .O(x60_y35),
    .I0(1'b0),
    .I1(x58_y38),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001110011010)
) lut_61_35 (
    .O(x61_y35),
    .I0(x59_y39),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101100000010)
) lut_62_35 (
    .O(x62_y35),
    .I0(x59_y37),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x60_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001100010011)
) lut_0_36 (
    .O(x0_y36),
    .I0(in1),
    .I1(in5),
    .I2(in8),
    .I3(in1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000100001000)
) lut_1_36 (
    .O(x1_y36),
    .I0(1'b0),
    .I1(in9),
    .I2(1'b0),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011000100001)
) lut_2_36 (
    .O(x2_y36),
    .I0(in7),
    .I1(1'b0),
    .I2(in4),
    .I3(in1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100011110100)
) lut_3_36 (
    .O(x3_y36),
    .I0(1'b0),
    .I1(in0),
    .I2(1'b0),
    .I3(in1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001110001111)
) lut_4_36 (
    .O(x4_y36),
    .I0(x2_y36),
    .I1(1'b0),
    .I2(x1_y35),
    .I3(x1_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110101000010)
) lut_5_36 (
    .O(x5_y36),
    .I0(x2_y31),
    .I1(1'b0),
    .I2(x3_y35),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011011000100)
) lut_6_36 (
    .O(x6_y36),
    .I0(x3_y41),
    .I1(x3_y32),
    .I2(1'b0),
    .I3(x4_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101011100011)
) lut_7_36 (
    .O(x7_y36),
    .I0(x5_y32),
    .I1(1'b0),
    .I2(x4_y34),
    .I3(x5_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011010100110)
) lut_8_36 (
    .O(x8_y36),
    .I0(x5_y37),
    .I1(x6_y40),
    .I2(x5_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110000000001)
) lut_9_36 (
    .O(x9_y36),
    .I0(x7_y41),
    .I1(1'b0),
    .I2(x5_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001001000001)
) lut_10_36 (
    .O(x10_y36),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x8_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110101110010)
) lut_11_36 (
    .O(x11_y36),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x8_y38),
    .I3(x8_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011011111101)
) lut_12_36 (
    .O(x12_y36),
    .I0(x10_y32),
    .I1(1'b0),
    .I2(x9_y33),
    .I3(x10_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000010111011)
) lut_13_36 (
    .O(x13_y36),
    .I0(1'b0),
    .I1(x10_y38),
    .I2(x11_y41),
    .I3(x11_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011100110011)
) lut_14_36 (
    .O(x14_y36),
    .I0(x11_y33),
    .I1(x11_y41),
    .I2(x11_y33),
    .I3(x11_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010011010010)
) lut_15_36 (
    .O(x15_y36),
    .I0(x13_y33),
    .I1(x13_y40),
    .I2(x12_y32),
    .I3(x13_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000101111010)
) lut_16_36 (
    .O(x16_y36),
    .I0(x13_y38),
    .I1(x13_y33),
    .I2(1'b0),
    .I3(x13_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101001010010)
) lut_17_36 (
    .O(x17_y36),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x14_y37),
    .I3(x14_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010100011010)
) lut_18_36 (
    .O(x18_y36),
    .I0(1'b0),
    .I1(x16_y38),
    .I2(x15_y38),
    .I3(x15_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101010110110)
) lut_19_36 (
    .O(x19_y36),
    .I0(x17_y33),
    .I1(x16_y36),
    .I2(x16_y34),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011010011100)
) lut_20_36 (
    .O(x20_y36),
    .I0(x17_y33),
    .I1(x18_y31),
    .I2(1'b0),
    .I3(x18_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101000001101)
) lut_21_36 (
    .O(x21_y36),
    .I0(x19_y32),
    .I1(x19_y38),
    .I2(1'b0),
    .I3(x19_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111011110011)
) lut_22_36 (
    .O(x22_y36),
    .I0(x20_y40),
    .I1(x20_y36),
    .I2(x20_y40),
    .I3(x20_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111100100000)
) lut_23_36 (
    .O(x23_y36),
    .I0(x20_y32),
    .I1(x20_y32),
    .I2(x21_y33),
    .I3(x21_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101000101001)
) lut_24_36 (
    .O(x24_y36),
    .I0(1'b0),
    .I1(x21_y40),
    .I2(x22_y36),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111111110010)
) lut_25_36 (
    .O(x25_y36),
    .I0(x23_y32),
    .I1(x22_y33),
    .I2(x23_y37),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010111100110)
) lut_26_36 (
    .O(x26_y36),
    .I0(x24_y31),
    .I1(x23_y40),
    .I2(x23_y40),
    .I3(x24_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101010101010)
) lut_27_36 (
    .O(x27_y36),
    .I0(x24_y36),
    .I1(x24_y35),
    .I2(x24_y41),
    .I3(x25_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000111011111)
) lut_28_36 (
    .O(x28_y36),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x25_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000100001110)
) lut_29_36 (
    .O(x29_y36),
    .I0(x26_y36),
    .I1(x27_y36),
    .I2(x26_y34),
    .I3(x26_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000000111101)
) lut_30_36 (
    .O(x30_y36),
    .I0(x27_y40),
    .I1(x27_y38),
    .I2(x27_y39),
    .I3(x27_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111111110011)
) lut_31_36 (
    .O(x31_y36),
    .I0(1'b0),
    .I1(x28_y39),
    .I2(x29_y31),
    .I3(x28_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110100000111)
) lut_32_36 (
    .O(x32_y36),
    .I0(1'b0),
    .I1(x30_y37),
    .I2(x29_y36),
    .I3(x29_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000110100011)
) lut_33_36 (
    .O(x33_y36),
    .I0(x30_y35),
    .I1(1'b0),
    .I2(x31_y36),
    .I3(x30_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111101100011)
) lut_34_36 (
    .O(x34_y36),
    .I0(x32_y31),
    .I1(x31_y33),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000000101000)
) lut_35_36 (
    .O(x35_y36),
    .I0(x32_y40),
    .I1(x32_y32),
    .I2(x33_y35),
    .I3(x33_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001010011000)
) lut_36_36 (
    .O(x36_y36),
    .I0(1'b0),
    .I1(x34_y38),
    .I2(1'b0),
    .I3(x33_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111100110111)
) lut_37_36 (
    .O(x37_y36),
    .I0(x35_y34),
    .I1(1'b0),
    .I2(x34_y37),
    .I3(x34_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000111110001)
) lut_38_36 (
    .O(x38_y36),
    .I0(x35_y40),
    .I1(x36_y37),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011111011100)
) lut_39_36 (
    .O(x39_y36),
    .I0(x36_y38),
    .I1(x37_y37),
    .I2(x36_y35),
    .I3(x36_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100110111100)
) lut_40_36 (
    .O(x40_y36),
    .I0(1'b0),
    .I1(x37_y31),
    .I2(1'b0),
    .I3(x38_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000000110111)
) lut_41_36 (
    .O(x41_y36),
    .I0(x39_y31),
    .I1(x39_y37),
    .I2(x38_y33),
    .I3(x38_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011000001101)
) lut_42_36 (
    .O(x42_y36),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x40_y35),
    .I3(x40_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010110010100)
) lut_43_36 (
    .O(x43_y36),
    .I0(x40_y35),
    .I1(x40_y40),
    .I2(x40_y38),
    .I3(x40_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111110101000)
) lut_44_36 (
    .O(x44_y36),
    .I0(x42_y36),
    .I1(x42_y33),
    .I2(x42_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110010110101)
) lut_45_36 (
    .O(x45_y36),
    .I0(x43_y33),
    .I1(x43_y32),
    .I2(x43_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111001111000)
) lut_46_36 (
    .O(x46_y36),
    .I0(x43_y35),
    .I1(x44_y40),
    .I2(1'b0),
    .I3(x43_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100011010101)
) lut_47_36 (
    .O(x47_y36),
    .I0(x44_y33),
    .I1(x44_y33),
    .I2(1'b0),
    .I3(x45_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000010000100)
) lut_48_36 (
    .O(x48_y36),
    .I0(x46_y37),
    .I1(x45_y33),
    .I2(x46_y35),
    .I3(x46_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110010000010)
) lut_49_36 (
    .O(x49_y36),
    .I0(x46_y39),
    .I1(x46_y38),
    .I2(x46_y33),
    .I3(x46_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000011101101)
) lut_50_36 (
    .O(x50_y36),
    .I0(x47_y40),
    .I1(x47_y32),
    .I2(x48_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001111010101)
) lut_51_36 (
    .O(x51_y36),
    .I0(x49_y38),
    .I1(x48_y41),
    .I2(x48_y37),
    .I3(x49_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110011110100)
) lut_52_36 (
    .O(x52_y36),
    .I0(x49_y35),
    .I1(x50_y37),
    .I2(x49_y32),
    .I3(x49_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100000011101)
) lut_53_36 (
    .O(x53_y36),
    .I0(x50_y38),
    .I1(x51_y39),
    .I2(x51_y41),
    .I3(x51_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110011000011)
) lut_54_36 (
    .O(x54_y36),
    .I0(x51_y39),
    .I1(x52_y32),
    .I2(x51_y39),
    .I3(x52_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010001111100)
) lut_55_36 (
    .O(x55_y36),
    .I0(x53_y40),
    .I1(x52_y34),
    .I2(x52_y39),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111000110110)
) lut_56_36 (
    .O(x56_y36),
    .I0(x54_y34),
    .I1(x54_y36),
    .I2(x54_y35),
    .I3(x54_y31)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010100110011)
) lut_57_36 (
    .O(x57_y36),
    .I0(x55_y32),
    .I1(x55_y34),
    .I2(x55_y33),
    .I3(x54_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011101101111)
) lut_58_36 (
    .O(x58_y36),
    .I0(x56_y40),
    .I1(x55_y31),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111110011110)
) lut_59_36 (
    .O(x59_y36),
    .I0(x56_y32),
    .I1(x57_y36),
    .I2(x56_y34),
    .I3(x56_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111010000111)
) lut_60_36 (
    .O(x60_y36),
    .I0(x57_y37),
    .I1(x58_y40),
    .I2(x57_y38),
    .I3(x57_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001110111000)
) lut_61_36 (
    .O(x61_y36),
    .I0(1'b0),
    .I1(x58_y38),
    .I2(1'b0),
    .I3(x59_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110100100100)
) lut_62_36 (
    .O(x62_y36),
    .I0(1'b0),
    .I1(x59_y39),
    .I2(1'b0),
    .I3(x60_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010011000011)
) lut_0_37 (
    .O(x0_y37),
    .I0(in4),
    .I1(in2),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111101001110)
) lut_1_37 (
    .O(x1_y37),
    .I0(in9),
    .I1(in7),
    .I2(in0),
    .I3(in5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100011101010)
) lut_2_37 (
    .O(x2_y37),
    .I0(in2),
    .I1(1'b0),
    .I2(1'b0),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110010101010)
) lut_3_37 (
    .O(x3_y37),
    .I0(in2),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110001101000)
) lut_4_37 (
    .O(x4_y37),
    .I0(x1_y33),
    .I1(x2_y39),
    .I2(x2_y33),
    .I3(x2_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000010101101)
) lut_5_37 (
    .O(x5_y37),
    .I0(1'b0),
    .I1(x2_y34),
    .I2(1'b0),
    .I3(x2_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101110100000)
) lut_6_37 (
    .O(x6_y37),
    .I0(1'b0),
    .I1(x3_y32),
    .I2(x4_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010100001110)
) lut_7_37 (
    .O(x7_y37),
    .I0(x4_y35),
    .I1(x4_y39),
    .I2(x4_y38),
    .I3(x4_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101001000001)
) lut_8_37 (
    .O(x8_y37),
    .I0(x5_y32),
    .I1(x6_y37),
    .I2(x5_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111000010001)
) lut_9_37 (
    .O(x9_y37),
    .I0(x7_y35),
    .I1(x7_y42),
    .I2(x5_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100101110110)
) lut_10_37 (
    .O(x10_y37),
    .I0(x8_y35),
    .I1(x8_y36),
    .I2(x8_y36),
    .I3(x7_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111011110111)
) lut_11_37 (
    .O(x11_y37),
    .I0(x8_y33),
    .I1(x8_y39),
    .I2(x9_y35),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111011010010)
) lut_12_37 (
    .O(x12_y37),
    .I0(x10_y42),
    .I1(x9_y40),
    .I2(1'b0),
    .I3(x10_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010000100101)
) lut_13_37 (
    .O(x13_y37),
    .I0(x11_y41),
    .I1(x11_y35),
    .I2(x10_y41),
    .I3(x11_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011001100001)
) lut_14_37 (
    .O(x14_y37),
    .I0(x12_y39),
    .I1(x12_y34),
    .I2(x12_y33),
    .I3(x11_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011110001111)
) lut_15_37 (
    .O(x15_y37),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x13_y41),
    .I3(x13_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000101011110)
) lut_16_37 (
    .O(x16_y37),
    .I0(x13_y32),
    .I1(x14_y33),
    .I2(x14_y33),
    .I3(x13_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010001101010)
) lut_17_37 (
    .O(x17_y37),
    .I0(x15_y42),
    .I1(x15_y35),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110010010100)
) lut_18_37 (
    .O(x18_y37),
    .I0(x15_y37),
    .I1(x16_y39),
    .I2(x16_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010010101100)
) lut_19_37 (
    .O(x19_y37),
    .I0(x16_y39),
    .I1(x17_y36),
    .I2(x16_y32),
    .I3(x17_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010011100101)
) lut_20_37 (
    .O(x20_y37),
    .I0(x18_y32),
    .I1(x17_y40),
    .I2(x17_y39),
    .I3(x17_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100101100011)
) lut_21_37 (
    .O(x21_y37),
    .I0(x18_y40),
    .I1(1'b0),
    .I2(x19_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010100100111)
) lut_22_37 (
    .O(x22_y37),
    .I0(1'b0),
    .I1(x20_y40),
    .I2(x20_y41),
    .I3(x20_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101100011110)
) lut_23_37 (
    .O(x23_y37),
    .I0(x20_y38),
    .I1(x21_y40),
    .I2(x20_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000110111110)
) lut_24_37 (
    .O(x24_y37),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x22_y38),
    .I3(x22_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110111110101)
) lut_25_37 (
    .O(x25_y37),
    .I0(1'b0),
    .I1(x23_y42),
    .I2(x23_y41),
    .I3(x22_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111001000100)
) lut_26_37 (
    .O(x26_y37),
    .I0(1'b0),
    .I1(x23_y38),
    .I2(x23_y38),
    .I3(x23_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111110101101)
) lut_27_37 (
    .O(x27_y37),
    .I0(x24_y38),
    .I1(x25_y34),
    .I2(1'b0),
    .I3(x25_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001111111010)
) lut_28_37 (
    .O(x28_y37),
    .I0(x25_y36),
    .I1(x25_y34),
    .I2(x25_y35),
    .I3(x26_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111111101010)
) lut_29_37 (
    .O(x29_y37),
    .I0(x26_y34),
    .I1(x27_y39),
    .I2(x27_y35),
    .I3(x27_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110100100110)
) lut_30_37 (
    .O(x30_y37),
    .I0(x28_y37),
    .I1(x28_y40),
    .I2(x28_y33),
    .I3(x27_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110010001010)
) lut_31_37 (
    .O(x31_y37),
    .I0(x29_y33),
    .I1(x28_y41),
    .I2(1'b0),
    .I3(x29_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111110010011)
) lut_32_37 (
    .O(x32_y37),
    .I0(x29_y33),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x30_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000011110100)
) lut_33_37 (
    .O(x33_y37),
    .I0(x30_y33),
    .I1(1'b0),
    .I2(x30_y38),
    .I3(x31_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011111111000)
) lut_34_37 (
    .O(x34_y37),
    .I0(x32_y39),
    .I1(1'b0),
    .I2(x32_y35),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011001000100)
) lut_35_37 (
    .O(x35_y37),
    .I0(x32_y38),
    .I1(x33_y35),
    .I2(x33_y40),
    .I3(x33_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000100001011)
) lut_36_37 (
    .O(x36_y37),
    .I0(1'b0),
    .I1(x33_y42),
    .I2(x33_y40),
    .I3(x33_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110101111111)
) lut_37_37 (
    .O(x37_y37),
    .I0(x35_y40),
    .I1(x34_y34),
    .I2(x35_y34),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010000000111)
) lut_38_37 (
    .O(x38_y37),
    .I0(x36_y41),
    .I1(x36_y36),
    .I2(1'b0),
    .I3(x35_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011010101010)
) lut_39_37 (
    .O(x39_y37),
    .I0(x36_y42),
    .I1(x36_y41),
    .I2(x36_y33),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001100010001)
) lut_40_37 (
    .O(x40_y37),
    .I0(x38_y37),
    .I1(x38_y42),
    .I2(x38_y38),
    .I3(x38_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110101101010)
) lut_41_37 (
    .O(x41_y37),
    .I0(x39_y42),
    .I1(x38_y39),
    .I2(x38_y35),
    .I3(x38_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100001110000)
) lut_42_37 (
    .O(x42_y37),
    .I0(x40_y35),
    .I1(x40_y36),
    .I2(1'b0),
    .I3(x39_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000111111000)
) lut_43_37 (
    .O(x43_y37),
    .I0(1'b0),
    .I1(x41_y39),
    .I2(x40_y36),
    .I3(x40_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111001101111)
) lut_44_37 (
    .O(x44_y37),
    .I0(1'b0),
    .I1(x41_y41),
    .I2(x41_y41),
    .I3(x42_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001111101010)
) lut_45_37 (
    .O(x45_y37),
    .I0(x43_y33),
    .I1(1'b0),
    .I2(x43_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001111110000)
) lut_46_37 (
    .O(x46_y37),
    .I0(x43_y32),
    .I1(x44_y36),
    .I2(1'b0),
    .I3(x43_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111000110100)
) lut_47_37 (
    .O(x47_y37),
    .I0(1'b0),
    .I1(x45_y42),
    .I2(x44_y32),
    .I3(x45_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000001010110)
) lut_48_37 (
    .O(x48_y37),
    .I0(x45_y40),
    .I1(x45_y36),
    .I2(1'b0),
    .I3(x46_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011110011101)
) lut_49_37 (
    .O(x49_y37),
    .I0(x46_y38),
    .I1(x46_y40),
    .I2(x47_y36),
    .I3(x46_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101000111000)
) lut_50_37 (
    .O(x50_y37),
    .I0(1'b0),
    .I1(x48_y32),
    .I2(x48_y37),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010110100011)
) lut_51_37 (
    .O(x51_y37),
    .I0(x49_y36),
    .I1(x48_y32),
    .I2(1'b0),
    .I3(x49_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101011100010)
) lut_52_37 (
    .O(x52_y37),
    .I0(x49_y32),
    .I1(1'b0),
    .I2(x49_y39),
    .I3(x50_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110101011001)
) lut_53_37 (
    .O(x53_y37),
    .I0(x50_y41),
    .I1(x51_y37),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101010001000)
) lut_54_37 (
    .O(x54_y37),
    .I0(x51_y34),
    .I1(x51_y33),
    .I2(x52_y40),
    .I3(x52_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010010011001)
) lut_55_37 (
    .O(x55_y37),
    .I0(1'b0),
    .I1(x53_y34),
    .I2(x52_y33),
    .I3(x52_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010011011000)
) lut_56_37 (
    .O(x56_y37),
    .I0(x53_y33),
    .I1(1'b0),
    .I2(x54_y36),
    .I3(x53_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011111010011)
) lut_57_37 (
    .O(x57_y37),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x55_y34),
    .I3(x55_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001101010100)
) lut_58_37 (
    .O(x58_y37),
    .I0(1'b0),
    .I1(x56_y37),
    .I2(x56_y37),
    .I3(x56_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011000110101)
) lut_59_37 (
    .O(x59_y37),
    .I0(x57_y39),
    .I1(x56_y39),
    .I2(x57_y41),
    .I3(x57_y32)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101000111100)
) lut_60_37 (
    .O(x60_y37),
    .I0(1'b0),
    .I1(x58_y37),
    .I2(x58_y33),
    .I3(x58_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110011101101)
) lut_61_37 (
    .O(x61_y37),
    .I0(x58_y33),
    .I1(x58_y37),
    .I2(x58_y37),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001011010001)
) lut_62_37 (
    .O(x62_y37),
    .I0(x60_y37),
    .I1(x60_y35),
    .I2(x59_y35),
    .I3(x60_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010001000111)
) lut_0_38 (
    .O(x0_y38),
    .I0(in0),
    .I1(in1),
    .I2(in0),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010010111001)
) lut_1_38 (
    .O(x1_y38),
    .I0(in1),
    .I1(in3),
    .I2(in0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010011000000)
) lut_2_38 (
    .O(x2_y38),
    .I0(1'b0),
    .I1(1'b0),
    .I2(in4),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011010001101)
) lut_3_38 (
    .O(x3_y38),
    .I0(in1),
    .I1(in6),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111101010100)
) lut_4_38 (
    .O(x4_y38),
    .I0(x2_y34),
    .I1(x1_y40),
    .I2(x1_y38),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110000010010)
) lut_5_38 (
    .O(x5_y38),
    .I0(x3_y34),
    .I1(x2_y36),
    .I2(x2_y41),
    .I3(x2_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110111110100)
) lut_6_38 (
    .O(x6_y38),
    .I0(1'b0),
    .I1(x4_y42),
    .I2(x3_y36),
    .I3(x3_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001010111110)
) lut_7_38 (
    .O(x7_y38),
    .I0(x5_y36),
    .I1(x5_y43),
    .I2(1'b0),
    .I3(x4_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100111000000)
) lut_8_38 (
    .O(x8_y38),
    .I0(x6_y42),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x5_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101110111011)
) lut_9_38 (
    .O(x9_y38),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x5_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011101101111)
) lut_10_38 (
    .O(x10_y38),
    .I0(x7_y38),
    .I1(x7_y40),
    .I2(1'b0),
    .I3(x7_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101000100110)
) lut_11_38 (
    .O(x11_y38),
    .I0(x9_y39),
    .I1(x9_y37),
    .I2(x8_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011001011011)
) lut_12_38 (
    .O(x12_y38),
    .I0(x10_y34),
    .I1(x9_y42),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010111100000)
) lut_13_38 (
    .O(x13_y38),
    .I0(x11_y37),
    .I1(1'b0),
    .I2(x10_y34),
    .I3(x10_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010010101110)
) lut_14_38 (
    .O(x14_y38),
    .I0(x12_y33),
    .I1(x12_y34),
    .I2(x12_y43),
    .I3(x12_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110001011000)
) lut_15_38 (
    .O(x15_y38),
    .I0(x13_y39),
    .I1(x12_y38),
    .I2(x13_y40),
    .I3(x13_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100000010011)
) lut_16_38 (
    .O(x16_y38),
    .I0(x14_y36),
    .I1(x13_y42),
    .I2(x14_y33),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101001101101)
) lut_17_38 (
    .O(x17_y38),
    .I0(x14_y43),
    .I1(x14_y39),
    .I2(x14_y37),
    .I3(x14_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000110110001)
) lut_18_38 (
    .O(x18_y38),
    .I0(x15_y39),
    .I1(x15_y33),
    .I2(x16_y34),
    .I3(x16_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010111011101)
) lut_19_38 (
    .O(x19_y38),
    .I0(1'b0),
    .I1(x17_y33),
    .I2(x17_y39),
    .I3(x16_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101111001001)
) lut_20_38 (
    .O(x20_y38),
    .I0(x17_y43),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111110110001)
) lut_21_38 (
    .O(x21_y38),
    .I0(x19_y42),
    .I1(x19_y35),
    .I2(x18_y36),
    .I3(x18_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100011011000)
) lut_22_38 (
    .O(x22_y38),
    .I0(1'b0),
    .I1(x19_y37),
    .I2(1'b0),
    .I3(x20_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010100111001)
) lut_23_38 (
    .O(x23_y38),
    .I0(x21_y33),
    .I1(x20_y33),
    .I2(x21_y34),
    .I3(x20_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000110101001)
) lut_24_38 (
    .O(x24_y38),
    .I0(x21_y33),
    .I1(x21_y41),
    .I2(x21_y34),
    .I3(x21_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010000001000)
) lut_25_38 (
    .O(x25_y38),
    .I0(x22_y38),
    .I1(1'b0),
    .I2(x22_y43),
    .I3(x23_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011000001010)
) lut_26_38 (
    .O(x26_y38),
    .I0(x24_y35),
    .I1(x24_y42),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011010001000)
) lut_27_38 (
    .O(x27_y38),
    .I0(x24_y43),
    .I1(x24_y36),
    .I2(x25_y34),
    .I3(x25_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010110010100)
) lut_28_38 (
    .O(x28_y38),
    .I0(x25_y34),
    .I1(x26_y38),
    .I2(x25_y39),
    .I3(x25_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100101100001)
) lut_29_38 (
    .O(x29_y38),
    .I0(x26_y40),
    .I1(x26_y33),
    .I2(x26_y39),
    .I3(x27_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001010000111)
) lut_30_38 (
    .O(x30_y38),
    .I0(x28_y43),
    .I1(x28_y34),
    .I2(x28_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100101101001)
) lut_31_38 (
    .O(x31_y38),
    .I0(x29_y36),
    .I1(x28_y39),
    .I2(x29_y42),
    .I3(x28_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111001000101)
) lut_32_38 (
    .O(x32_y38),
    .I0(x29_y35),
    .I1(x29_y33),
    .I2(x29_y41),
    .I3(x29_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010000001111)
) lut_33_38 (
    .O(x33_y38),
    .I0(x30_y42),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x30_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110010101011)
) lut_34_38 (
    .O(x34_y38),
    .I0(x31_y33),
    .I1(x32_y34),
    .I2(1'b0),
    .I3(x32_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001101010100)
) lut_35_38 (
    .O(x35_y38),
    .I0(x33_y38),
    .I1(1'b0),
    .I2(x33_y34),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101101100010)
) lut_36_38 (
    .O(x36_y38),
    .I0(x34_y33),
    .I1(x34_y33),
    .I2(x34_y42),
    .I3(x33_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001011111101)
) lut_37_38 (
    .O(x37_y38),
    .I0(x35_y41),
    .I1(x35_y42),
    .I2(1'b0),
    .I3(x35_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111111011001)
) lut_38_38 (
    .O(x38_y38),
    .I0(x35_y37),
    .I1(x36_y41),
    .I2(x36_y35),
    .I3(x35_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110000001101)
) lut_39_38 (
    .O(x39_y38),
    .I0(x36_y34),
    .I1(x36_y40),
    .I2(1'b0),
    .I3(x36_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110110010101)
) lut_40_38 (
    .O(x40_y38),
    .I0(x38_y42),
    .I1(x38_y38),
    .I2(x37_y36),
    .I3(x37_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100000000000)
) lut_41_38 (
    .O(x41_y38),
    .I0(x38_y39),
    .I1(1'b0),
    .I2(x39_y38),
    .I3(x39_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001100001001)
) lut_42_38 (
    .O(x42_y38),
    .I0(x39_y41),
    .I1(x39_y42),
    .I2(x40_y33),
    .I3(x39_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100001011001)
) lut_43_38 (
    .O(x43_y38),
    .I0(x40_y38),
    .I1(x40_y33),
    .I2(x40_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011110010110)
) lut_44_38 (
    .O(x44_y38),
    .I0(1'b0),
    .I1(x42_y33),
    .I2(x42_y42),
    .I3(x42_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010100100011)
) lut_45_38 (
    .O(x45_y38),
    .I0(x42_y39),
    .I1(1'b0),
    .I2(x42_y36),
    .I3(x42_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001001001011)
) lut_46_38 (
    .O(x46_y38),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x43_y35),
    .I3(x44_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111010110000)
) lut_47_38 (
    .O(x47_y38),
    .I0(x44_y33),
    .I1(x45_y35),
    .I2(1'b0),
    .I3(x44_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111010100011)
) lut_48_38 (
    .O(x48_y38),
    .I0(1'b0),
    .I1(x46_y37),
    .I2(x45_y36),
    .I3(x45_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001111100011)
) lut_49_38 (
    .O(x49_y38),
    .I0(1'b0),
    .I1(x46_y39),
    .I2(1'b0),
    .I3(x46_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110010001000)
) lut_50_38 (
    .O(x50_y38),
    .I0(x48_y37),
    .I1(x47_y36),
    .I2(x48_y38),
    .I3(x48_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100010001011)
) lut_51_38 (
    .O(x51_y38),
    .I0(x49_y34),
    .I1(1'b0),
    .I2(x48_y42),
    .I3(x49_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000011100101)
) lut_52_38 (
    .O(x52_y38),
    .I0(1'b0),
    .I1(x49_y40),
    .I2(x49_y38),
    .I3(x49_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000011001101)
) lut_53_38 (
    .O(x53_y38),
    .I0(x50_y33),
    .I1(x50_y36),
    .I2(x50_y41),
    .I3(x50_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101110110010)
) lut_54_38 (
    .O(x54_y38),
    .I0(x51_y42),
    .I1(x51_y42),
    .I2(x52_y33),
    .I3(x52_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000100110101)
) lut_55_38 (
    .O(x55_y38),
    .I0(x53_y42),
    .I1(x53_y42),
    .I2(x52_y42),
    .I3(x53_y33)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110001110010)
) lut_56_38 (
    .O(x56_y38),
    .I0(x53_y41),
    .I1(1'b0),
    .I2(x54_y43),
    .I3(x53_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011100011110)
) lut_57_38 (
    .O(x57_y38),
    .I0(x54_y37),
    .I1(x54_y39),
    .I2(x54_y38),
    .I3(x55_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010011111100)
) lut_58_38 (
    .O(x58_y38),
    .I0(x55_y36),
    .I1(x55_y37),
    .I2(1'b0),
    .I3(x56_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000101100101)
) lut_59_38 (
    .O(x59_y38),
    .I0(x56_y37),
    .I1(x57_y37),
    .I2(x56_y41),
    .I3(x57_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011101110000)
) lut_60_38 (
    .O(x60_y38),
    .I0(x58_y43),
    .I1(x57_y41),
    .I2(x57_y34),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101100001011)
) lut_61_38 (
    .O(x61_y38),
    .I0(1'b0),
    .I1(x59_y41),
    .I2(x59_y38),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000100011011)
) lut_62_38 (
    .O(x62_y38),
    .I0(x59_y34),
    .I1(x60_y36),
    .I2(x60_y41),
    .I3(x60_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001010010101)
) lut_0_39 (
    .O(x0_y39),
    .I0(in3),
    .I1(1'b0),
    .I2(in4),
    .I3(in9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111011011101)
) lut_1_39 (
    .O(x1_y39),
    .I0(in2),
    .I1(in9),
    .I2(in2),
    .I3(in3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011011001010)
) lut_2_39 (
    .O(x2_y39),
    .I0(in0),
    .I1(in4),
    .I2(in1),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100110110001)
) lut_3_39 (
    .O(x3_y39),
    .I0(in7),
    .I1(1'b0),
    .I2(x1_y37),
    .I3(in5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101110100110)
) lut_4_39 (
    .O(x4_y39),
    .I0(1'b0),
    .I1(x2_y35),
    .I2(1'b0),
    .I3(x1_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011111110101)
) lut_5_39 (
    .O(x5_y39),
    .I0(x3_y43),
    .I1(x3_y44),
    .I2(x3_y41),
    .I3(x2_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011000100100)
) lut_6_39 (
    .O(x6_y39),
    .I0(x3_y34),
    .I1(x3_y43),
    .I2(x3_y39),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110001011011)
) lut_7_39 (
    .O(x7_y39),
    .I0(x5_y39),
    .I1(x4_y43),
    .I2(x4_y36),
    .I3(x4_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110011110100)
) lut_8_39 (
    .O(x8_y39),
    .I0(1'b0),
    .I1(x6_y42),
    .I2(x6_y39),
    .I3(x5_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111110101010)
) lut_9_39 (
    .O(x9_y39),
    .I0(x6_y39),
    .I1(x6_y34),
    .I2(x6_y39),
    .I3(x5_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011111111101)
) lut_10_39 (
    .O(x10_y39),
    .I0(x7_y38),
    .I1(1'b0),
    .I2(x8_y43),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100001100110)
) lut_11_39 (
    .O(x11_y39),
    .I0(x9_y44),
    .I1(x9_y41),
    .I2(x8_y41),
    .I3(x8_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110010110110)
) lut_12_39 (
    .O(x12_y39),
    .I0(x10_y43),
    .I1(x10_y43),
    .I2(x10_y43),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111100001011)
) lut_13_39 (
    .O(x13_y39),
    .I0(x11_y40),
    .I1(x10_y42),
    .I2(x11_y40),
    .I3(x11_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110101111110)
) lut_14_39 (
    .O(x14_y39),
    .I0(1'b0),
    .I1(x11_y38),
    .I2(1'b0),
    .I3(x12_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001111101100)
) lut_15_39 (
    .O(x15_y39),
    .I0(x13_y39),
    .I1(x12_y38),
    .I2(x13_y43),
    .I3(x12_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011110111101)
) lut_16_39 (
    .O(x16_y39),
    .I0(x14_y35),
    .I1(x14_y38),
    .I2(x14_y41),
    .I3(x14_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011101001010)
) lut_17_39 (
    .O(x17_y39),
    .I0(x14_y34),
    .I1(x14_y35),
    .I2(x14_y40),
    .I3(x14_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111100110000)
) lut_18_39 (
    .O(x18_y39),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x16_y39),
    .I3(x16_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000000011001)
) lut_19_39 (
    .O(x19_y39),
    .I0(x17_y41),
    .I1(x17_y43),
    .I2(1'b0),
    .I3(x16_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010010001111)
) lut_20_39 (
    .O(x20_y39),
    .I0(x18_y36),
    .I1(x17_y39),
    .I2(x17_y42),
    .I3(x18_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101111001110)
) lut_21_39 (
    .O(x21_y39),
    .I0(x18_y40),
    .I1(x18_y39),
    .I2(1'b0),
    .I3(x19_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101000000101)
) lut_22_39 (
    .O(x22_y39),
    .I0(x19_y44),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x20_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100110100010)
) lut_23_39 (
    .O(x23_y39),
    .I0(1'b0),
    .I1(x21_y42),
    .I2(x21_y38),
    .I3(x21_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101000101110)
) lut_24_39 (
    .O(x24_y39),
    .I0(x22_y41),
    .I1(x21_y38),
    .I2(1'b0),
    .I3(x22_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001110000100)
) lut_25_39 (
    .O(x25_y39),
    .I0(1'b0),
    .I1(x23_y43),
    .I2(x22_y42),
    .I3(x23_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110111100101)
) lut_26_39 (
    .O(x26_y39),
    .I0(x24_y38),
    .I1(x24_y41),
    .I2(x24_y36),
    .I3(x24_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110111000111)
) lut_27_39 (
    .O(x27_y39),
    .I0(x24_y36),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x24_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010100111111)
) lut_28_39 (
    .O(x28_y39),
    .I0(1'b0),
    .I1(x26_y39),
    .I2(x26_y44),
    .I3(x25_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110001110001)
) lut_29_39 (
    .O(x29_y39),
    .I0(x26_y37),
    .I1(x26_y42),
    .I2(x26_y36),
    .I3(x26_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110000010101)
) lut_30_39 (
    .O(x30_y39),
    .I0(1'b0),
    .I1(x27_y36),
    .I2(x28_y39),
    .I3(x27_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101001111000)
) lut_31_39 (
    .O(x31_y39),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x28_y40),
    .I3(x29_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111110001101)
) lut_32_39 (
    .O(x32_y39),
    .I0(x29_y38),
    .I1(x29_y41),
    .I2(x29_y38),
    .I3(x30_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011001000010)
) lut_33_39 (
    .O(x33_y39),
    .I0(1'b0),
    .I1(x30_y43),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111101001001)
) lut_34_39 (
    .O(x34_y39),
    .I0(x32_y44),
    .I1(1'b0),
    .I2(x31_y43),
    .I3(x32_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010000110111)
) lut_35_39 (
    .O(x35_y39),
    .I0(x33_y44),
    .I1(x33_y42),
    .I2(x32_y35),
    .I3(x33_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000000011100)
) lut_36_39 (
    .O(x36_y39),
    .I0(x34_y39),
    .I1(x33_y40),
    .I2(x34_y44),
    .I3(x34_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000010100011)
) lut_37_39 (
    .O(x37_y39),
    .I0(x34_y37),
    .I1(x35_y44),
    .I2(x35_y37),
    .I3(x34_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010000110011)
) lut_38_39 (
    .O(x38_y39),
    .I0(1'b0),
    .I1(x36_y34),
    .I2(x35_y36),
    .I3(x35_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011000001100)
) lut_39_39 (
    .O(x39_y39),
    .I0(x36_y41),
    .I1(x37_y43),
    .I2(x37_y42),
    .I3(x36_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000100000101)
) lut_40_39 (
    .O(x40_y39),
    .I0(x37_y35),
    .I1(1'b0),
    .I2(x37_y37),
    .I3(x38_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001001011111)
) lut_41_39 (
    .O(x41_y39),
    .I0(1'b0),
    .I1(x39_y41),
    .I2(x39_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000000001010)
) lut_42_39 (
    .O(x42_y39),
    .I0(x40_y42),
    .I1(x39_y42),
    .I2(1'b0),
    .I3(x40_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101101101100)
) lut_43_39 (
    .O(x43_y39),
    .I0(x40_y41),
    .I1(1'b0),
    .I2(x41_y36),
    .I3(x40_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110011011110)
) lut_44_39 (
    .O(x44_y39),
    .I0(x42_y44),
    .I1(x41_y38),
    .I2(1'b0),
    .I3(x42_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101110000110)
) lut_45_39 (
    .O(x45_y39),
    .I0(x43_y43),
    .I1(x42_y41),
    .I2(x43_y37),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110100100000)
) lut_46_39 (
    .O(x46_y39),
    .I0(1'b0),
    .I1(x44_y41),
    .I2(x43_y38),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001100110001)
) lut_47_39 (
    .O(x47_y39),
    .I0(1'b0),
    .I1(x44_y34),
    .I2(x45_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011001001100)
) lut_48_39 (
    .O(x48_y39),
    .I0(x45_y42),
    .I1(x46_y41),
    .I2(x46_y41),
    .I3(x45_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100101111110)
) lut_49_39 (
    .O(x49_y39),
    .I0(x46_y39),
    .I1(x46_y37),
    .I2(x46_y34),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111101010010)
) lut_50_39 (
    .O(x50_y39),
    .I0(1'b0),
    .I1(x48_y36),
    .I2(x48_y37),
    .I3(x48_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110110011010)
) lut_51_39 (
    .O(x51_y39),
    .I0(x49_y41),
    .I1(x49_y35),
    .I2(1'b0),
    .I3(x49_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010010110011)
) lut_52_39 (
    .O(x52_y39),
    .I0(x49_y44),
    .I1(x49_y42),
    .I2(x49_y37),
    .I3(x50_y34)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100001101111)
) lut_53_39 (
    .O(x53_y39),
    .I0(x50_y41),
    .I1(1'b0),
    .I2(x50_y36),
    .I3(x51_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111110101101)
) lut_54_39 (
    .O(x54_y39),
    .I0(x52_y40),
    .I1(x51_y37),
    .I2(x52_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100001100011)
) lut_55_39 (
    .O(x55_y39),
    .I0(1'b0),
    .I1(x53_y39),
    .I2(x52_y43),
    .I3(x52_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101111101001)
) lut_56_39 (
    .O(x56_y39),
    .I0(x54_y34),
    .I1(x53_y43),
    .I2(x53_y37),
    .I3(x54_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100010011001)
) lut_57_39 (
    .O(x57_y39),
    .I0(x55_y39),
    .I1(x54_y44),
    .I2(x54_y40),
    .I3(x54_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100010010001)
) lut_58_39 (
    .O(x58_y39),
    .I0(x56_y35),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x56_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010111111111)
) lut_59_39 (
    .O(x59_y39),
    .I0(x57_y37),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010000110111)
) lut_60_39 (
    .O(x60_y39),
    .I0(x58_y41),
    .I1(x57_y39),
    .I2(1'b0),
    .I3(x57_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000101110011)
) lut_61_39 (
    .O(x61_y39),
    .I0(x59_y43),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x58_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000000101001)
) lut_62_39 (
    .O(x62_y39),
    .I0(x59_y44),
    .I1(x60_y41),
    .I2(x59_y40),
    .I3(x60_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001111000011)
) lut_0_40 (
    .O(x0_y40),
    .I0(in1),
    .I1(in5),
    .I2(in8),
    .I3(in9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000101001101)
) lut_1_40 (
    .O(x1_y40),
    .I0(1'b0),
    .I1(in3),
    .I2(in0),
    .I3(in5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111111101000)
) lut_2_40 (
    .O(x2_y40),
    .I0(in6),
    .I1(in8),
    .I2(in4),
    .I3(in6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000110010001)
) lut_3_40 (
    .O(x3_y40),
    .I0(in9),
    .I1(in6),
    .I2(in3),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111000011111)
) lut_4_40 (
    .O(x4_y40),
    .I0(x2_y36),
    .I1(x1_y40),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010110010010)
) lut_5_40 (
    .O(x5_y40),
    .I0(x3_y37),
    .I1(x3_y38),
    .I2(x2_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111101000011)
) lut_6_40 (
    .O(x6_y40),
    .I0(1'b0),
    .I1(x3_y41),
    .I2(x3_y36),
    .I3(x3_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110111011110)
) lut_7_40 (
    .O(x7_y40),
    .I0(1'b0),
    .I1(x4_y37),
    .I2(x4_y37),
    .I3(x5_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001110010111)
) lut_8_40 (
    .O(x8_y40),
    .I0(x6_y45),
    .I1(x5_y35),
    .I2(1'b0),
    .I3(x5_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100111001000)
) lut_9_40 (
    .O(x9_y40),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x5_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111101100100)
) lut_10_40 (
    .O(x10_y40),
    .I0(x8_y40),
    .I1(x8_y44),
    .I2(x7_y35),
    .I3(x7_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100110001001)
) lut_11_40 (
    .O(x11_y40),
    .I0(x8_y42),
    .I1(x9_y42),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011100011110)
) lut_12_40 (
    .O(x12_y40),
    .I0(1'b0),
    .I1(x10_y38),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011101100011)
) lut_13_40 (
    .O(x13_y40),
    .I0(x11_y41),
    .I1(x10_y35),
    .I2(1'b0),
    .I3(x10_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001011100010)
) lut_14_40 (
    .O(x14_y40),
    .I0(x12_y39),
    .I1(x11_y43),
    .I2(x11_y38),
    .I3(x12_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011111011100)
) lut_15_40 (
    .O(x15_y40),
    .I0(x12_y44),
    .I1(x13_y41),
    .I2(x13_y39),
    .I3(x12_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001000001111)
) lut_16_40 (
    .O(x16_y40),
    .I0(x14_y35),
    .I1(x13_y37),
    .I2(1'b0),
    .I3(x13_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001001011010)
) lut_17_40 (
    .O(x17_y40),
    .I0(x15_y44),
    .I1(x14_y37),
    .I2(x15_y41),
    .I3(x14_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101011001111)
) lut_18_40 (
    .O(x18_y40),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x16_y40),
    .I3(x16_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011011110110)
) lut_19_40 (
    .O(x19_y40),
    .I0(1'b0),
    .I1(x17_y39),
    .I2(x17_y38),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101100101011)
) lut_20_40 (
    .O(x20_y40),
    .I0(x17_y45),
    .I1(x17_y38),
    .I2(x18_y36),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001010100001)
) lut_21_40 (
    .O(x21_y40),
    .I0(1'b0),
    .I1(x19_y37),
    .I2(x18_y38),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100000100100)
) lut_22_40 (
    .O(x22_y40),
    .I0(x19_y42),
    .I1(x19_y35),
    .I2(x19_y42),
    .I3(x19_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111011101001)
) lut_23_40 (
    .O(x23_y40),
    .I0(1'b0),
    .I1(x20_y40),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110101111111)
) lut_24_40 (
    .O(x24_y40),
    .I0(x22_y42),
    .I1(x22_y39),
    .I2(1'b0),
    .I3(x21_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110011000100)
) lut_25_40 (
    .O(x25_y40),
    .I0(x23_y38),
    .I1(1'b0),
    .I2(x22_y37),
    .I3(x22_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100001010101)
) lut_26_40 (
    .O(x26_y40),
    .I0(x24_y35),
    .I1(x24_y37),
    .I2(x24_y40),
    .I3(x24_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101110100001)
) lut_27_40 (
    .O(x27_y40),
    .I0(x24_y41),
    .I1(x25_y44),
    .I2(x25_y45),
    .I3(x25_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001110110001)
) lut_28_40 (
    .O(x28_y40),
    .I0(x26_y37),
    .I1(x25_y44),
    .I2(x26_y44),
    .I3(x25_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000011111000)
) lut_29_40 (
    .O(x29_y40),
    .I0(1'b0),
    .I1(x27_y40),
    .I2(x26_y36),
    .I3(x26_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110010001000)
) lut_30_40 (
    .O(x30_y40),
    .I0(1'b0),
    .I1(x28_y40),
    .I2(x27_y44),
    .I3(x27_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000101101110)
) lut_31_40 (
    .O(x31_y40),
    .I0(x29_y43),
    .I1(x28_y41),
    .I2(x29_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010011101001)
) lut_32_40 (
    .O(x32_y40),
    .I0(x29_y40),
    .I1(x29_y45),
    .I2(x29_y45),
    .I3(x30_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001111110011)
) lut_33_40 (
    .O(x33_y40),
    .I0(x30_y40),
    .I1(x31_y43),
    .I2(x30_y39),
    .I3(x30_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010100101010)
) lut_34_40 (
    .O(x34_y40),
    .I0(x31_y42),
    .I1(x32_y35),
    .I2(x32_y44),
    .I3(x32_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111101010111)
) lut_35_40 (
    .O(x35_y40),
    .I0(x32_y42),
    .I1(x32_y37),
    .I2(x33_y35),
    .I3(x32_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101111010111)
) lut_36_40 (
    .O(x36_y40),
    .I0(x34_y41),
    .I1(x34_y39),
    .I2(x34_y45),
    .I3(x33_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000100110010)
) lut_37_40 (
    .O(x37_y40),
    .I0(x34_y39),
    .I1(x34_y37),
    .I2(x35_y44),
    .I3(x34_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010010110000)
) lut_38_40 (
    .O(x38_y40),
    .I0(x36_y39),
    .I1(x36_y44),
    .I2(x36_y40),
    .I3(x36_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100011011101)
) lut_39_40 (
    .O(x39_y40),
    .I0(x36_y38),
    .I1(x37_y40),
    .I2(x36_y44),
    .I3(x36_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011111001111)
) lut_40_40 (
    .O(x40_y40),
    .I0(x38_y37),
    .I1(1'b0),
    .I2(x38_y43),
    .I3(x38_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110001010101)
) lut_41_40 (
    .O(x41_y40),
    .I0(x39_y36),
    .I1(1'b0),
    .I2(x39_y41),
    .I3(x38_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101010011001)
) lut_42_40 (
    .O(x42_y40),
    .I0(x39_y35),
    .I1(x39_y44),
    .I2(x39_y44),
    .I3(x39_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111101001100)
) lut_43_40 (
    .O(x43_y40),
    .I0(x40_y37),
    .I1(1'b0),
    .I2(x41_y39),
    .I3(x40_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111111000110)
) lut_44_40 (
    .O(x44_y40),
    .I0(x41_y42),
    .I1(x42_y43),
    .I2(x41_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111101110100)
) lut_45_40 (
    .O(x45_y40),
    .I0(x43_y40),
    .I1(x42_y42),
    .I2(x42_y37),
    .I3(x42_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110101100111)
) lut_46_40 (
    .O(x46_y40),
    .I0(1'b0),
    .I1(x44_y42),
    .I2(x44_y43),
    .I3(x43_y35)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011001000011)
) lut_47_40 (
    .O(x47_y40),
    .I0(x45_y35),
    .I1(x45_y39),
    .I2(1'b0),
    .I3(x44_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011111011110)
) lut_48_40 (
    .O(x48_y40),
    .I0(x45_y43),
    .I1(1'b0),
    .I2(x45_y45),
    .I3(x45_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100010101001)
) lut_49_40 (
    .O(x49_y40),
    .I0(x46_y43),
    .I1(x47_y36),
    .I2(x46_y39),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101110100101)
) lut_50_40 (
    .O(x50_y40),
    .I0(1'b0),
    .I1(x47_y43),
    .I2(x48_y35),
    .I3(x47_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010010001000)
) lut_51_40 (
    .O(x51_y40),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x48_y39),
    .I3(x48_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111001110111)
) lut_52_40 (
    .O(x52_y40),
    .I0(1'b0),
    .I1(x50_y41),
    .I2(x50_y35),
    .I3(x49_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111100001110)
) lut_53_40 (
    .O(x53_y40),
    .I0(x51_y39),
    .I1(x50_y36),
    .I2(x50_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011101010010)
) lut_54_40 (
    .O(x54_y40),
    .I0(1'b0),
    .I1(x52_y38),
    .I2(x51_y36),
    .I3(x51_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111000110011)
) lut_55_40 (
    .O(x55_y40),
    .I0(x52_y42),
    .I1(x53_y42),
    .I2(1'b0),
    .I3(x52_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001100110111)
) lut_56_40 (
    .O(x56_y40),
    .I0(x54_y35),
    .I1(x53_y36),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110110100010)
) lut_57_40 (
    .O(x57_y40),
    .I0(x55_y45),
    .I1(x54_y36),
    .I2(x55_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010100011010)
) lut_58_40 (
    .O(x58_y40),
    .I0(x56_y40),
    .I1(x55_y40),
    .I2(x56_y36),
    .I3(x55_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101110110001)
) lut_59_40 (
    .O(x59_y40),
    .I0(1'b0),
    .I1(x57_y45),
    .I2(1'b0),
    .I3(x56_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001110110010)
) lut_60_40 (
    .O(x60_y40),
    .I0(1'b0),
    .I1(x57_y44),
    .I2(x58_y36),
    .I3(x58_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101110001110)
) lut_61_40 (
    .O(x61_y40),
    .I0(x58_y35),
    .I1(x59_y38),
    .I2(x58_y37),
    .I3(x59_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011011001100)
) lut_62_40 (
    .O(x62_y40),
    .I0(x60_y39),
    .I1(x59_y36),
    .I2(x59_y42),
    .I3(x60_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001101110001)
) lut_0_41 (
    .O(x0_y41),
    .I0(in2),
    .I1(in4),
    .I2(in0),
    .I3(in4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111001010001)
) lut_1_41 (
    .O(x1_y41),
    .I0(in3),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100010000100)
) lut_2_41 (
    .O(x2_y41),
    .I0(in4),
    .I1(in3),
    .I2(1'b0),
    .I3(in1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001101010001)
) lut_3_41 (
    .O(x3_y41),
    .I0(in5),
    .I1(1'b0),
    .I2(in6),
    .I3(x1_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001001000000)
) lut_4_41 (
    .O(x4_y41),
    .I0(x1_y44),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010010000100)
) lut_5_41 (
    .O(x5_y41),
    .I0(1'b0),
    .I1(x2_y43),
    .I2(1'b0),
    .I3(x3_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011000010001)
) lut_6_41 (
    .O(x6_y41),
    .I0(x4_y40),
    .I1(x3_y43),
    .I2(1'b0),
    .I3(x3_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101110100100)
) lut_7_41 (
    .O(x7_y41),
    .I0(x5_y46),
    .I1(x4_y40),
    .I2(1'b0),
    .I3(x5_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100000101010)
) lut_8_41 (
    .O(x8_y41),
    .I0(x5_y37),
    .I1(x5_y39),
    .I2(x6_y43),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011000011000)
) lut_9_41 (
    .O(x9_y41),
    .I0(x6_y42),
    .I1(x7_y44),
    .I2(x6_y43),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110111100001)
) lut_10_41 (
    .O(x10_y41),
    .I0(x7_y46),
    .I1(x7_y43),
    .I2(x7_y41),
    .I3(x8_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011101001111)
) lut_11_41 (
    .O(x11_y41),
    .I0(x9_y45),
    .I1(1'b0),
    .I2(x8_y46),
    .I3(x8_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000100011110)
) lut_12_41 (
    .O(x12_y41),
    .I0(x9_y46),
    .I1(x10_y39),
    .I2(x9_y45),
    .I3(x10_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000010111111)
) lut_13_41 (
    .O(x13_y41),
    .I0(x11_y41),
    .I1(1'b0),
    .I2(x11_y36),
    .I3(x11_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110010001110)
) lut_14_41 (
    .O(x14_y41),
    .I0(x12_y43),
    .I1(x11_y39),
    .I2(1'b0),
    .I3(x11_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110100110010)
) lut_15_41 (
    .O(x15_y41),
    .I0(x12_y36),
    .I1(x13_y44),
    .I2(x13_y41),
    .I3(x12_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100011101101)
) lut_16_41 (
    .O(x16_y41),
    .I0(1'b0),
    .I1(x13_y43),
    .I2(x13_y39),
    .I3(x13_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111000001010)
) lut_17_41 (
    .O(x17_y41),
    .I0(x14_y38),
    .I1(x14_y42),
    .I2(x15_y41),
    .I3(x15_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111011101111)
) lut_18_41 (
    .O(x18_y41),
    .I0(x15_y46),
    .I1(1'b0),
    .I2(x16_y41),
    .I3(x15_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011100000000)
) lut_19_41 (
    .O(x19_y41),
    .I0(x17_y40),
    .I1(x17_y45),
    .I2(x16_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111101000100)
) lut_20_41 (
    .O(x20_y41),
    .I0(x17_y38),
    .I1(1'b0),
    .I2(x18_y36),
    .I3(x17_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010110010000)
) lut_21_41 (
    .O(x21_y41),
    .I0(1'b0),
    .I1(x18_y45),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011011111001)
) lut_22_41 (
    .O(x22_y41),
    .I0(x19_y46),
    .I1(x19_y45),
    .I2(x19_y38),
    .I3(x19_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111101010010)
) lut_23_41 (
    .O(x23_y41),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x20_y39),
    .I3(x20_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101110100000)
) lut_24_41 (
    .O(x24_y41),
    .I0(1'b0),
    .I1(x22_y38),
    .I2(x22_y44),
    .I3(x21_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111111110111)
) lut_25_41 (
    .O(x25_y41),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x22_y36),
    .I3(x23_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010100001000)
) lut_26_41 (
    .O(x26_y41),
    .I0(x24_y38),
    .I1(x24_y38),
    .I2(x23_y37),
    .I3(x24_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101101001110)
) lut_27_41 (
    .O(x27_y41),
    .I0(x25_y37),
    .I1(x24_y46),
    .I2(x25_y41),
    .I3(x24_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101111101101)
) lut_28_41 (
    .O(x28_y41),
    .I0(1'b0),
    .I1(x26_y43),
    .I2(x25_y42),
    .I3(x26_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111011110111)
) lut_29_41 (
    .O(x29_y41),
    .I0(x27_y39),
    .I1(x26_y44),
    .I2(x26_y44),
    .I3(x27_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000010110011)
) lut_30_41 (
    .O(x30_y41),
    .I0(x28_y36),
    .I1(x28_y42),
    .I2(1'b0),
    .I3(x27_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000011100011)
) lut_31_41 (
    .O(x31_y41),
    .I0(x29_y36),
    .I1(x28_y43),
    .I2(x28_y38),
    .I3(x28_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010001001110)
) lut_32_41 (
    .O(x32_y41),
    .I0(x29_y43),
    .I1(x30_y42),
    .I2(x29_y46),
    .I3(x29_y36)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011100011001)
) lut_33_41 (
    .O(x33_y41),
    .I0(x30_y42),
    .I1(x31_y43),
    .I2(x31_y39),
    .I3(x31_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010001001110)
) lut_34_41 (
    .O(x34_y41),
    .I0(x31_y40),
    .I1(x31_y38),
    .I2(x31_y39),
    .I3(x31_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010111000111)
) lut_35_41 (
    .O(x35_y41),
    .I0(x32_y38),
    .I1(1'b0),
    .I2(x33_y44),
    .I3(x32_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101110000011)
) lut_36_41 (
    .O(x36_y41),
    .I0(1'b0),
    .I1(x34_y45),
    .I2(x33_y38),
    .I3(x34_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010111100001)
) lut_37_41 (
    .O(x37_y41),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x34_y39),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111100000100)
) lut_38_41 (
    .O(x38_y41),
    .I0(1'b0),
    .I1(x35_y37),
    .I2(1'b0),
    .I3(x35_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111011010001)
) lut_39_41 (
    .O(x39_y41),
    .I0(1'b0),
    .I1(x36_y44),
    .I2(x36_y37),
    .I3(x36_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011110110111)
) lut_40_41 (
    .O(x40_y41),
    .I0(1'b0),
    .I1(x38_y42),
    .I2(x37_y38),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011100100101)
) lut_41_41 (
    .O(x41_y41),
    .I0(x39_y46),
    .I1(x38_y40),
    .I2(x39_y39),
    .I3(x39_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011110011000)
) lut_42_41 (
    .O(x42_y41),
    .I0(x39_y37),
    .I1(x40_y44),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101101101010)
) lut_43_41 (
    .O(x43_y41),
    .I0(x40_y38),
    .I1(1'b0),
    .I2(x40_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001010110100)
) lut_44_41 (
    .O(x44_y41),
    .I0(x42_y45),
    .I1(1'b0),
    .I2(x42_y36),
    .I3(x42_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110101111100)
) lut_45_41 (
    .O(x45_y41),
    .I0(x43_y44),
    .I1(x43_y39),
    .I2(x43_y40),
    .I3(x42_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000010010111)
) lut_46_41 (
    .O(x46_y41),
    .I0(x43_y39),
    .I1(x44_y40),
    .I2(1'b0),
    .I3(x43_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100000100110)
) lut_47_41 (
    .O(x47_y41),
    .I0(x45_y36),
    .I1(x44_y44),
    .I2(x44_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010101111010)
) lut_48_41 (
    .O(x48_y41),
    .I0(x46_y38),
    .I1(x46_y43),
    .I2(x46_y38),
    .I3(x45_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001111000001)
) lut_49_41 (
    .O(x49_y41),
    .I0(1'b0),
    .I1(x46_y46),
    .I2(x47_y43),
    .I3(x47_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110000010100)
) lut_50_41 (
    .O(x50_y41),
    .I0(x48_y36),
    .I1(x47_y39),
    .I2(x48_y39),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110011010111)
) lut_51_41 (
    .O(x51_y41),
    .I0(x49_y40),
    .I1(x48_y42),
    .I2(1'b0),
    .I3(x48_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010010010001)
) lut_52_41 (
    .O(x52_y41),
    .I0(x49_y42),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x50_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001111010010)
) lut_53_41 (
    .O(x53_y41),
    .I0(1'b0),
    .I1(x50_y42),
    .I2(x50_y38),
    .I3(x50_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001000101111)
) lut_54_41 (
    .O(x54_y41),
    .I0(x52_y44),
    .I1(x51_y38),
    .I2(x51_y40),
    .I3(x52_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111110101000)
) lut_55_41 (
    .O(x55_y41),
    .I0(x53_y41),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x53_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010011111000)
) lut_56_41 (
    .O(x56_y41),
    .I0(1'b0),
    .I1(x54_y42),
    .I2(x53_y40),
    .I3(x54_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011100011000)
) lut_57_41 (
    .O(x57_y41),
    .I0(x55_y43),
    .I1(x55_y38),
    .I2(x54_y41),
    .I3(x54_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101110000001)
) lut_58_41 (
    .O(x58_y41),
    .I0(x56_y46),
    .I1(x56_y41),
    .I2(x55_y45),
    .I3(x56_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101111010111)
) lut_59_41 (
    .O(x59_y41),
    .I0(x57_y37),
    .I1(x57_y41),
    .I2(x56_y40),
    .I3(x57_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110010100000)
) lut_60_41 (
    .O(x60_y41),
    .I0(x57_y38),
    .I1(x57_y39),
    .I2(x58_y46),
    .I3(x58_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001111111111)
) lut_61_41 (
    .O(x61_y41),
    .I0(x58_y44),
    .I1(x59_y38),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011111100100)
) lut_62_41 (
    .O(x62_y41),
    .I0(1'b0),
    .I1(x60_y43),
    .I2(1'b0),
    .I3(x59_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011100101001)
) lut_0_42 (
    .O(x0_y42),
    .I0(1'b0),
    .I1(in6),
    .I2(in6),
    .I3(in6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101000100011)
) lut_1_42 (
    .O(x1_y42),
    .I0(in7),
    .I1(1'b0),
    .I2(in3),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001001001000)
) lut_2_42 (
    .O(x2_y42),
    .I0(in0),
    .I1(in6),
    .I2(in2),
    .I3(in7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100110000010)
) lut_3_42 (
    .O(x3_y42),
    .I0(in3),
    .I1(1'b0),
    .I2(in9),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110100111011)
) lut_4_42 (
    .O(x4_y42),
    .I0(x2_y45),
    .I1(x1_y47),
    .I2(x2_y44),
    .I3(x1_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100000011110)
) lut_5_42 (
    .O(x5_y42),
    .I0(x2_y37),
    .I1(x2_y38),
    .I2(x3_y45),
    .I3(x2_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000001110010)
) lut_6_42 (
    .O(x6_y42),
    .I0(x4_y46),
    .I1(x3_y38),
    .I2(1'b0),
    .I3(x4_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001101101110)
) lut_7_42 (
    .O(x7_y42),
    .I0(x4_y47),
    .I1(x4_y47),
    .I2(x5_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100101011111)
) lut_8_42 (
    .O(x8_y42),
    .I0(x6_y41),
    .I1(1'b0),
    .I2(x6_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101111110000)
) lut_9_42 (
    .O(x9_y42),
    .I0(1'b0),
    .I1(x6_y45),
    .I2(x6_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101100001110)
) lut_10_42 (
    .O(x10_y42),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x7_y47),
    .I3(x8_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011011011100)
) lut_11_42 (
    .O(x11_y42),
    .I0(x9_y38),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x8_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001100101000)
) lut_12_42 (
    .O(x12_y42),
    .I0(x10_y45),
    .I1(x10_y46),
    .I2(x10_y43),
    .I3(x9_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110000110001)
) lut_13_42 (
    .O(x13_y42),
    .I0(x11_y46),
    .I1(x10_y42),
    .I2(x11_y42),
    .I3(x11_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011101001101)
) lut_14_42 (
    .O(x14_y42),
    .I0(x12_y39),
    .I1(x11_y43),
    .I2(x12_y38),
    .I3(x12_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011001011100)
) lut_15_42 (
    .O(x15_y42),
    .I0(x13_y46),
    .I1(x12_y42),
    .I2(1'b0),
    .I3(x12_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111111111111)
) lut_16_42 (
    .O(x16_y42),
    .I0(x14_y40),
    .I1(x14_y37),
    .I2(x13_y45),
    .I3(x14_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111001111000)
) lut_17_42 (
    .O(x17_y42),
    .I0(x15_y47),
    .I1(x15_y44),
    .I2(1'b0),
    .I3(x14_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010111110010)
) lut_18_42 (
    .O(x18_y42),
    .I0(x16_y37),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111111000110)
) lut_19_42 (
    .O(x19_y42),
    .I0(x17_y39),
    .I1(x16_y38),
    .I2(x16_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101011001000)
) lut_20_42 (
    .O(x20_y42),
    .I0(x18_y46),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001011011010)
) lut_21_42 (
    .O(x21_y42),
    .I0(x18_y47),
    .I1(x19_y41),
    .I2(x18_y46),
    .I3(x19_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011100011010)
) lut_22_42 (
    .O(x22_y42),
    .I0(x20_y40),
    .I1(1'b0),
    .I2(x20_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101011001000)
) lut_23_42 (
    .O(x23_y42),
    .I0(x20_y45),
    .I1(1'b0),
    .I2(x20_y47),
    .I3(x21_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001101001010)
) lut_24_42 (
    .O(x24_y42),
    .I0(x22_y37),
    .I1(1'b0),
    .I2(x22_y45),
    .I3(x22_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011011001111)
) lut_25_42 (
    .O(x25_y42),
    .I0(x22_y37),
    .I1(x23_y44),
    .I2(1'b0),
    .I3(x23_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011101001000)
) lut_26_42 (
    .O(x26_y42),
    .I0(x24_y39),
    .I1(x24_y41),
    .I2(1'b0),
    .I3(x24_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000101011110)
) lut_27_42 (
    .O(x27_y42),
    .I0(x24_y43),
    .I1(x24_y47),
    .I2(1'b0),
    .I3(x24_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100011010011)
) lut_28_42 (
    .O(x28_y42),
    .I0(x26_y38),
    .I1(1'b0),
    .I2(x26_y47),
    .I3(x26_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010000101101)
) lut_29_42 (
    .O(x29_y42),
    .I0(x26_y39),
    .I1(1'b0),
    .I2(x26_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011110110010)
) lut_30_42 (
    .O(x30_y42),
    .I0(x28_y45),
    .I1(x27_y37),
    .I2(x28_y43),
    .I3(x28_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111001010100)
) lut_31_42 (
    .O(x31_y42),
    .I0(x28_y39),
    .I1(x29_y43),
    .I2(x29_y43),
    .I3(x28_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110010001000)
) lut_32_42 (
    .O(x32_y42),
    .I0(x30_y37),
    .I1(x29_y43),
    .I2(1'b0),
    .I3(x30_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111010000100)
) lut_33_42 (
    .O(x33_y42),
    .I0(x30_y39),
    .I1(x30_y39),
    .I2(x31_y43),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110101101110)
) lut_34_42 (
    .O(x34_y42),
    .I0(x32_y39),
    .I1(x32_y38),
    .I2(x32_y38),
    .I3(x31_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011111011111)
) lut_35_42 (
    .O(x35_y42),
    .I0(x32_y38),
    .I1(x32_y40),
    .I2(x32_y38),
    .I3(x32_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000111101001)
) lut_36_42 (
    .O(x36_y42),
    .I0(x33_y41),
    .I1(x34_y39),
    .I2(x34_y40),
    .I3(x33_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011010000100)
) lut_37_42 (
    .O(x37_y42),
    .I0(x34_y46),
    .I1(x34_y38),
    .I2(1'b0),
    .I3(x34_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101110110011)
) lut_38_42 (
    .O(x38_y42),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000111111011)
) lut_39_42 (
    .O(x39_y42),
    .I0(x37_y43),
    .I1(x37_y43),
    .I2(x37_y41),
    .I3(x37_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001111110110)
) lut_40_42 (
    .O(x40_y42),
    .I0(1'b0),
    .I1(x38_y42),
    .I2(x37_y45),
    .I3(x38_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000111100010)
) lut_41_42 (
    .O(x41_y42),
    .I0(x38_y38),
    .I1(x39_y41),
    .I2(x38_y37),
    .I3(x38_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010001011001)
) lut_42_42 (
    .O(x42_y42),
    .I0(1'b0),
    .I1(x39_y37),
    .I2(x40_y46),
    .I3(x39_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110001111001)
) lut_43_42 (
    .O(x43_y42),
    .I0(x40_y46),
    .I1(1'b0),
    .I2(x41_y47),
    .I3(x40_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001110010001)
) lut_44_42 (
    .O(x44_y42),
    .I0(x42_y42),
    .I1(1'b0),
    .I2(x41_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000011001110)
) lut_45_42 (
    .O(x45_y42),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x42_y40),
    .I3(x42_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000010110001)
) lut_46_42 (
    .O(x46_y42),
    .I0(x43_y38),
    .I1(x43_y42),
    .I2(1'b0),
    .I3(x43_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110010100111)
) lut_47_42 (
    .O(x47_y42),
    .I0(x44_y45),
    .I1(x45_y40),
    .I2(1'b0),
    .I3(x44_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010000010101)
) lut_48_42 (
    .O(x48_y42),
    .I0(1'b0),
    .I1(x45_y41),
    .I2(x45_y43),
    .I3(x46_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100111110000)
) lut_49_42 (
    .O(x49_y42),
    .I0(x46_y47),
    .I1(x47_y47),
    .I2(1'b0),
    .I3(x47_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110011111110)
) lut_50_42 (
    .O(x50_y42),
    .I0(x47_y44),
    .I1(x47_y39),
    .I2(x47_y46),
    .I3(x47_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101101101101)
) lut_51_42 (
    .O(x51_y42),
    .I0(x48_y46),
    .I1(x49_y37),
    .I2(x48_y47),
    .I3(x49_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101100100110)
) lut_52_42 (
    .O(x52_y42),
    .I0(x50_y44),
    .I1(x49_y42),
    .I2(x49_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110100100100)
) lut_53_42 (
    .O(x53_y42),
    .I0(1'b0),
    .I1(x50_y40),
    .I2(x51_y38),
    .I3(x51_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000101000110)
) lut_54_42 (
    .O(x54_y42),
    .I0(x51_y38),
    .I1(x52_y38),
    .I2(x51_y37),
    .I3(x51_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100100001111)
) lut_55_42 (
    .O(x55_y42),
    .I0(1'b0),
    .I1(x53_y40),
    .I2(x53_y38),
    .I3(x53_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101001111101)
) lut_56_42 (
    .O(x56_y42),
    .I0(x54_y46),
    .I1(x53_y38),
    .I2(x54_y45),
    .I3(x54_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011001010111)
) lut_57_42 (
    .O(x57_y42),
    .I0(x54_y37),
    .I1(x54_y39),
    .I2(x55_y47),
    .I3(x55_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000101101100)
) lut_58_42 (
    .O(x58_y42),
    .I0(1'b0),
    .I1(x55_y40),
    .I2(x56_y40),
    .I3(x56_y37)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000011011111)
) lut_59_42 (
    .O(x59_y42),
    .I0(x57_y38),
    .I1(x56_y41),
    .I2(1'b0),
    .I3(x57_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101111110001)
) lut_60_42 (
    .O(x60_y42),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x57_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110001011111)
) lut_61_42 (
    .O(x61_y42),
    .I0(x59_y42),
    .I1(x59_y38),
    .I2(x59_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011101000011)
) lut_62_42 (
    .O(x62_y42),
    .I0(x59_y39),
    .I1(1'b0),
    .I2(x59_y40),
    .I3(x59_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000111000111)
) lut_0_43 (
    .O(x0_y43),
    .I0(in3),
    .I1(1'b0),
    .I2(in2),
    .I3(in5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000011110011)
) lut_1_43 (
    .O(x1_y43),
    .I0(1'b0),
    .I1(in5),
    .I2(1'b0),
    .I3(in4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010010110000)
) lut_2_43 (
    .O(x2_y43),
    .I0(in9),
    .I1(1'b0),
    .I2(in9),
    .I3(in7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000011100100)
) lut_3_43 (
    .O(x3_y43),
    .I0(x1_y46),
    .I1(1'b0),
    .I2(x1_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111001010001)
) lut_4_43 (
    .O(x4_y43),
    .I0(x2_y48),
    .I1(x1_y48),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100000011000)
) lut_5_43 (
    .O(x5_y43),
    .I0(1'b0),
    .I1(x3_y47),
    .I2(1'b0),
    .I3(x3_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010000010101)
) lut_6_43 (
    .O(x6_y43),
    .I0(1'b0),
    .I1(x3_y47),
    .I2(x4_y47),
    .I3(x3_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111000101010)
) lut_7_43 (
    .O(x7_y43),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x5_y44),
    .I3(x4_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111000100111)
) lut_8_43 (
    .O(x8_y43),
    .I0(x5_y44),
    .I1(1'b0),
    .I2(x6_y41),
    .I3(x5_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100100001011)
) lut_9_43 (
    .O(x9_y43),
    .I0(x7_y38),
    .I1(x7_y48),
    .I2(x6_y41),
    .I3(x5_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000100011100)
) lut_10_43 (
    .O(x10_y43),
    .I0(x8_y47),
    .I1(1'b0),
    .I2(x8_y40),
    .I3(x8_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100011000111)
) lut_11_43 (
    .O(x11_y43),
    .I0(x8_y39),
    .I1(x8_y41),
    .I2(x9_y45),
    .I3(x8_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010010001011)
) lut_12_43 (
    .O(x12_y43),
    .I0(x9_y44),
    .I1(x10_y42),
    .I2(x9_y39),
    .I3(x9_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100001010011)
) lut_13_43 (
    .O(x13_y43),
    .I0(x10_y39),
    .I1(x10_y42),
    .I2(x10_y46),
    .I3(x11_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010001000000)
) lut_14_43 (
    .O(x14_y43),
    .I0(x12_y43),
    .I1(x12_y43),
    .I2(x12_y40),
    .I3(x12_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100111011101)
) lut_15_43 (
    .O(x15_y43),
    .I0(x13_y47),
    .I1(x13_y42),
    .I2(x13_y39),
    .I3(x12_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001100011100)
) lut_16_43 (
    .O(x16_y43),
    .I0(x13_y40),
    .I1(x13_y48),
    .I2(x13_y41),
    .I3(x13_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010110011100)
) lut_17_43 (
    .O(x17_y43),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x15_y48),
    .I3(x15_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000110111110)
) lut_18_43 (
    .O(x18_y43),
    .I0(x16_y48),
    .I1(x15_y40),
    .I2(1'b0),
    .I3(x16_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000101001011)
) lut_19_43 (
    .O(x19_y43),
    .I0(x16_y39),
    .I1(x16_y38),
    .I2(x16_y38),
    .I3(x17_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010100011111)
) lut_20_43 (
    .O(x20_y43),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x17_y44),
    .I3(x18_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000101011001)
) lut_21_43 (
    .O(x21_y43),
    .I0(x18_y41),
    .I1(x19_y40),
    .I2(x18_y40),
    .I3(x18_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101101000110)
) lut_22_43 (
    .O(x22_y43),
    .I0(x20_y48),
    .I1(x19_y48),
    .I2(1'b0),
    .I3(x19_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001100110111)
) lut_23_43 (
    .O(x23_y43),
    .I0(x21_y46),
    .I1(x20_y46),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010000101001)
) lut_24_43 (
    .O(x24_y43),
    .I0(x21_y48),
    .I1(x22_y48),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110010111101)
) lut_25_43 (
    .O(x25_y43),
    .I0(x23_y48),
    .I1(x22_y38),
    .I2(x23_y43),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100010100110)
) lut_26_43 (
    .O(x26_y43),
    .I0(x24_y41),
    .I1(x23_y42),
    .I2(x23_y48),
    .I3(x24_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000011111100)
) lut_27_43 (
    .O(x27_y43),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110111111000)
) lut_28_43 (
    .O(x28_y43),
    .I0(x25_y48),
    .I1(x25_y44),
    .I2(x25_y38),
    .I3(x25_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111111001010)
) lut_29_43 (
    .O(x29_y43),
    .I0(x27_y41),
    .I1(1'b0),
    .I2(x27_y46),
    .I3(x27_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011100000111)
) lut_30_43 (
    .O(x30_y43),
    .I0(x27_y44),
    .I1(1'b0),
    .I2(x28_y46),
    .I3(x28_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001010110110)
) lut_31_43 (
    .O(x31_y43),
    .I0(1'b0),
    .I1(x29_y39),
    .I2(1'b0),
    .I3(x28_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100110001101)
) lut_32_43 (
    .O(x32_y43),
    .I0(x29_y45),
    .I1(x29_y43),
    .I2(x29_y46),
    .I3(x29_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000111111110)
) lut_33_43 (
    .O(x33_y43),
    .I0(1'b0),
    .I1(x31_y38),
    .I2(x31_y46),
    .I3(x31_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110101000000)
) lut_34_43 (
    .O(x34_y43),
    .I0(x32_y44),
    .I1(x32_y40),
    .I2(1'b0),
    .I3(x32_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111011001011)
) lut_35_43 (
    .O(x35_y43),
    .I0(x32_y44),
    .I1(x32_y42),
    .I2(x33_y48),
    .I3(x32_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001011110001)
) lut_36_43 (
    .O(x36_y43),
    .I0(x33_y42),
    .I1(x33_y48),
    .I2(1'b0),
    .I3(x33_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010010001010)
) lut_37_43 (
    .O(x37_y43),
    .I0(x34_y39),
    .I1(x35_y47),
    .I2(x35_y41),
    .I3(x35_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011100101110)
) lut_38_43 (
    .O(x38_y43),
    .I0(x36_y38),
    .I1(1'b0),
    .I2(x35_y42),
    .I3(x36_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100001101000)
) lut_39_43 (
    .O(x39_y43),
    .I0(x37_y40),
    .I1(x37_y45),
    .I2(x37_y40),
    .I3(x37_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110111001001)
) lut_40_43 (
    .O(x40_y43),
    .I0(x38_y42),
    .I1(x38_y38),
    .I2(x38_y44),
    .I3(x37_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110101000001)
) lut_41_43 (
    .O(x41_y43),
    .I0(x39_y40),
    .I1(x39_y42),
    .I2(x39_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110101010000)
) lut_42_43 (
    .O(x42_y43),
    .I0(x39_y43),
    .I1(x40_y47),
    .I2(x39_y41),
    .I3(x39_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110101111110)
) lut_43_43 (
    .O(x43_y43),
    .I0(1'b0),
    .I1(x41_y48),
    .I2(x40_y44),
    .I3(x41_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101001111111)
) lut_44_43 (
    .O(x44_y43),
    .I0(x42_y42),
    .I1(x41_y47),
    .I2(x41_y38),
    .I3(x41_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000011111010)
) lut_45_43 (
    .O(x45_y43),
    .I0(x43_y44),
    .I1(x43_y48),
    .I2(x42_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110110011101)
) lut_46_43 (
    .O(x46_y43),
    .I0(x43_y43),
    .I1(x43_y45),
    .I2(1'b0),
    .I3(x43_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010010101011)
) lut_47_43 (
    .O(x47_y43),
    .I0(x44_y46),
    .I1(1'b0),
    .I2(x44_y39),
    .I3(x44_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110001110001)
) lut_48_43 (
    .O(x48_y43),
    .I0(x46_y41),
    .I1(x46_y45),
    .I2(x45_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101101001010)
) lut_49_43 (
    .O(x49_y43),
    .I0(x47_y40),
    .I1(x46_y39),
    .I2(x47_y40),
    .I3(x47_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111101000010)
) lut_50_43 (
    .O(x50_y43),
    .I0(x47_y48),
    .I1(1'b0),
    .I2(x48_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110010001111)
) lut_51_43 (
    .O(x51_y43),
    .I0(1'b0),
    .I1(x49_y43),
    .I2(x49_y47),
    .I3(x48_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100110011101)
) lut_52_43 (
    .O(x52_y43),
    .I0(x49_y46),
    .I1(x49_y40),
    .I2(1'b0),
    .I3(x50_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100101000001)
) lut_53_43 (
    .O(x53_y43),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x50_y45),
    .I3(x51_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100111100101)
) lut_54_43 (
    .O(x54_y43),
    .I0(x51_y43),
    .I1(x52_y42),
    .I2(x52_y46),
    .I3(x51_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010000111001)
) lut_55_43 (
    .O(x55_y43),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x53_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000100011111)
) lut_56_43 (
    .O(x56_y43),
    .I0(x53_y45),
    .I1(1'b0),
    .I2(x54_y42),
    .I3(x53_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001011100100)
) lut_57_43 (
    .O(x57_y43),
    .I0(1'b0),
    .I1(x55_y43),
    .I2(x55_y42),
    .I3(x54_y38)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011110111110)
) lut_58_43 (
    .O(x58_y43),
    .I0(1'b0),
    .I1(x55_y40),
    .I2(1'b0),
    .I3(x55_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100000100101)
) lut_59_43 (
    .O(x59_y43),
    .I0(x57_y45),
    .I1(x57_y45),
    .I2(x57_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100100111101)
) lut_60_43 (
    .O(x60_y43),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x57_y41),
    .I3(x58_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100011110110)
) lut_61_43 (
    .O(x61_y43),
    .I0(x58_y41),
    .I1(x58_y38),
    .I2(x59_y40),
    .I3(x58_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011101101100)
) lut_62_43 (
    .O(x62_y43),
    .I0(x59_y44),
    .I1(x60_y39),
    .I2(1'b0),
    .I3(x59_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010100110100)
) lut_0_44 (
    .O(x0_y44),
    .I0(in0),
    .I1(in9),
    .I2(in9),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010110100100)
) lut_1_44 (
    .O(x1_y44),
    .I0(1'b0),
    .I1(1'b0),
    .I2(in9),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101000101000)
) lut_2_44 (
    .O(x2_y44),
    .I0(in2),
    .I1(in6),
    .I2(in0),
    .I3(in9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100000111010)
) lut_3_44 (
    .O(x3_y44),
    .I0(x1_y46),
    .I1(in3),
    .I2(in6),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101110111111)
) lut_4_44 (
    .O(x4_y44),
    .I0(x2_y40),
    .I1(1'b0),
    .I2(x1_y45),
    .I3(x2_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011011110001)
) lut_5_44 (
    .O(x5_y44),
    .I0(1'b0),
    .I1(x2_y49),
    .I2(x2_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000111110101)
) lut_6_44 (
    .O(x6_y44),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x3_y48),
    .I3(x4_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000000001110)
) lut_7_44 (
    .O(x7_y44),
    .I0(x4_y43),
    .I1(x4_y44),
    .I2(x4_y47),
    .I3(x5_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010011100111)
) lut_8_44 (
    .O(x8_y44),
    .I0(x6_y45),
    .I1(x5_y49),
    .I2(x5_y46),
    .I3(x5_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000010010000)
) lut_9_44 (
    .O(x9_y44),
    .I0(x6_y49),
    .I1(x7_y49),
    .I2(x5_y46),
    .I3(x5_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111001011000)
) lut_10_44 (
    .O(x10_y44),
    .I0(x8_y39),
    .I1(x7_y48),
    .I2(1'b0),
    .I3(x7_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011110000001)
) lut_11_44 (
    .O(x11_y44),
    .I0(x9_y46),
    .I1(1'b0),
    .I2(x9_y47),
    .I3(x9_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100110000111)
) lut_12_44 (
    .O(x12_y44),
    .I0(x9_y39),
    .I1(x10_y49),
    .I2(x10_y48),
    .I3(x9_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000101100011)
) lut_13_44 (
    .O(x13_y44),
    .I0(x11_y44),
    .I1(1'b0),
    .I2(x10_y40),
    .I3(x10_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010001100110)
) lut_14_44 (
    .O(x14_y44),
    .I0(x12_y41),
    .I1(1'b0),
    .I2(x11_y39),
    .I3(x12_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010100001000)
) lut_15_44 (
    .O(x15_y44),
    .I0(x13_y42),
    .I1(x13_y46),
    .I2(x12_y40),
    .I3(x13_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000010011010)
) lut_16_44 (
    .O(x16_y44),
    .I0(x13_y47),
    .I1(x13_y41),
    .I2(x13_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111011010100)
) lut_17_44 (
    .O(x17_y44),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x15_y47),
    .I3(x14_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101001111011)
) lut_18_44 (
    .O(x18_y44),
    .I0(1'b0),
    .I1(x15_y40),
    .I2(x16_y47),
    .I3(x15_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111100100010)
) lut_19_44 (
    .O(x19_y44),
    .I0(x16_y49),
    .I1(x17_y48),
    .I2(x17_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001101110100)
) lut_20_44 (
    .O(x20_y44),
    .I0(x17_y43),
    .I1(x17_y42),
    .I2(x18_y46),
    .I3(x17_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011100111100)
) lut_21_44 (
    .O(x21_y44),
    .I0(1'b0),
    .I1(x19_y44),
    .I2(x19_y46),
    .I3(x18_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011000101100)
) lut_22_44 (
    .O(x22_y44),
    .I0(1'b0),
    .I1(x19_y45),
    .I2(1'b0),
    .I3(x19_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010101000000)
) lut_23_44 (
    .O(x23_y44),
    .I0(x21_y41),
    .I1(x21_y39),
    .I2(x21_y44),
    .I3(x21_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111011001001)
) lut_24_44 (
    .O(x24_y44),
    .I0(x22_y41),
    .I1(x21_y46),
    .I2(x21_y47),
    .I3(x21_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000100010101)
) lut_25_44 (
    .O(x25_y44),
    .I0(1'b0),
    .I1(x22_y42),
    .I2(x22_y44),
    .I3(x23_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010110011000)
) lut_26_44 (
    .O(x26_y44),
    .I0(x24_y40),
    .I1(1'b0),
    .I2(x24_y41),
    .I3(x24_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001100000111)
) lut_27_44 (
    .O(x27_y44),
    .I0(x25_y48),
    .I1(x25_y49),
    .I2(x24_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001011100111)
) lut_28_44 (
    .O(x28_y44),
    .I0(1'b0),
    .I1(x26_y41),
    .I2(x25_y48),
    .I3(x26_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011100101001)
) lut_29_44 (
    .O(x29_y44),
    .I0(x27_y48),
    .I1(x27_y40),
    .I2(x27_y39),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100110111001)
) lut_30_44 (
    .O(x30_y44),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011000101001)
) lut_31_44 (
    .O(x31_y44),
    .I0(1'b0),
    .I1(x28_y40),
    .I2(x28_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101000110100)
) lut_32_44 (
    .O(x32_y44),
    .I0(x29_y48),
    .I1(x30_y44),
    .I2(x30_y44),
    .I3(x30_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110010100100)
) lut_33_44 (
    .O(x33_y44),
    .I0(x30_y48),
    .I1(x30_y41),
    .I2(x31_y49),
    .I3(x31_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000110100110)
) lut_34_44 (
    .O(x34_y44),
    .I0(1'b0),
    .I1(x31_y47),
    .I2(x31_y46),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110010101111)
) lut_35_44 (
    .O(x35_y44),
    .I0(1'b0),
    .I1(x32_y43),
    .I2(x33_y39),
    .I3(x32_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110000110000)
) lut_36_44 (
    .O(x36_y44),
    .I0(1'b0),
    .I1(x33_y47),
    .I2(x33_y44),
    .I3(x33_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111001101000)
) lut_37_44 (
    .O(x37_y44),
    .I0(x35_y43),
    .I1(x35_y44),
    .I2(x34_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010111000110)
) lut_38_44 (
    .O(x38_y44),
    .I0(x36_y41),
    .I1(x36_y44),
    .I2(x36_y44),
    .I3(x35_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010011010011)
) lut_39_44 (
    .O(x39_y44),
    .I0(x36_y46),
    .I1(x37_y40),
    .I2(x36_y46),
    .I3(x36_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011101100000)
) lut_40_44 (
    .O(x40_y44),
    .I0(x38_y42),
    .I1(x38_y42),
    .I2(1'b0),
    .I3(x38_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101111001101)
) lut_41_44 (
    .O(x41_y44),
    .I0(x39_y49),
    .I1(x39_y44),
    .I2(1'b0),
    .I3(x39_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010010110101)
) lut_42_44 (
    .O(x42_y44),
    .I0(x40_y43),
    .I1(x39_y45),
    .I2(x39_y40),
    .I3(x40_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100110110010)
) lut_43_44 (
    .O(x43_y44),
    .I0(x41_y40),
    .I1(1'b0),
    .I2(x41_y49),
    .I3(x40_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000000110100)
) lut_44_44 (
    .O(x44_y44),
    .I0(x41_y45),
    .I1(x41_y45),
    .I2(1'b0),
    .I3(x41_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011100010001)
) lut_45_44 (
    .O(x45_y44),
    .I0(x43_y41),
    .I1(1'b0),
    .I2(x43_y39),
    .I3(x42_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001010001001)
) lut_46_44 (
    .O(x46_y44),
    .I0(x43_y39),
    .I1(x43_y41),
    .I2(x44_y47),
    .I3(x44_y40)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000101000000)
) lut_47_44 (
    .O(x47_y44),
    .I0(x45_y45),
    .I1(x45_y40),
    .I2(1'b0),
    .I3(x44_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101111010110)
) lut_48_44 (
    .O(x48_y44),
    .I0(x45_y39),
    .I1(x46_y40),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110000001101)
) lut_49_44 (
    .O(x49_y44),
    .I0(x46_y44),
    .I1(x47_y44),
    .I2(x47_y47),
    .I3(x47_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110011010000)
) lut_50_44 (
    .O(x50_y44),
    .I0(x48_y46),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x47_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111101011010)
) lut_51_44 (
    .O(x51_y44),
    .I0(1'b0),
    .I1(x48_y44),
    .I2(x49_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010010000011)
) lut_52_44 (
    .O(x52_y44),
    .I0(x50_y44),
    .I1(x50_y47),
    .I2(x50_y48),
    .I3(x49_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011000100100)
) lut_53_44 (
    .O(x53_y44),
    .I0(x50_y48),
    .I1(1'b0),
    .I2(x51_y46),
    .I3(x51_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010010000011)
) lut_54_44 (
    .O(x54_y44),
    .I0(1'b0),
    .I1(x51_y43),
    .I2(1'b0),
    .I3(x51_y39)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010000010011)
) lut_55_44 (
    .O(x55_y44),
    .I0(1'b0),
    .I1(x53_y44),
    .I2(x53_y47),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011111000001)
) lut_56_44 (
    .O(x56_y44),
    .I0(x54_y44),
    .I1(1'b0),
    .I2(x54_y43),
    .I3(x54_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111100101001)
) lut_57_44 (
    .O(x57_y44),
    .I0(1'b0),
    .I1(x55_y40),
    .I2(x55_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110010001111)
) lut_58_44 (
    .O(x58_y44),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x55_y49),
    .I3(x56_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010000101100)
) lut_59_44 (
    .O(x59_y44),
    .I0(x56_y39),
    .I1(x56_y40),
    .I2(x57_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001001111110)
) lut_60_44 (
    .O(x60_y44),
    .I0(x57_y45),
    .I1(1'b0),
    .I2(x58_y49),
    .I3(x58_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000111001000)
) lut_61_44 (
    .O(x61_y44),
    .I0(x59_y39),
    .I1(1'b0),
    .I2(x59_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010000011001)
) lut_62_44 (
    .O(x62_y44),
    .I0(x59_y45),
    .I1(x60_y40),
    .I2(x60_y39),
    .I3(x59_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010101101011)
) lut_0_45 (
    .O(x0_y45),
    .I0(in0),
    .I1(1'b0),
    .I2(in1),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100011011010)
) lut_1_45 (
    .O(x1_y45),
    .I0(in6),
    .I1(in2),
    .I2(1'b0),
    .I3(in3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101100111011)
) lut_2_45 (
    .O(x2_y45),
    .I0(in1),
    .I1(1'b0),
    .I2(in1),
    .I3(in6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101000010010)
) lut_3_45 (
    .O(x3_y45),
    .I0(in4),
    .I1(x1_y47),
    .I2(1'b0),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100011111111)
) lut_4_45 (
    .O(x4_y45),
    .I0(x1_y47),
    .I1(x2_y47),
    .I2(x2_y45),
    .I3(x2_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010000101101)
) lut_5_45 (
    .O(x5_y45),
    .I0(x3_y42),
    .I1(x3_y43),
    .I2(x2_y47),
    .I3(x3_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101110110010)
) lut_6_45 (
    .O(x6_y45),
    .I0(x4_y47),
    .I1(x3_y45),
    .I2(x3_y43),
    .I3(x3_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001110101111)
) lut_7_45 (
    .O(x7_y45),
    .I0(x4_y48),
    .I1(x4_y48),
    .I2(x4_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001101111000)
) lut_8_45 (
    .O(x8_y45),
    .I0(1'b0),
    .I1(x6_y50),
    .I2(x5_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010110101010)
) lut_9_45 (
    .O(x9_y45),
    .I0(x6_y40),
    .I1(1'b0),
    .I2(x5_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111011010011)
) lut_10_45 (
    .O(x10_y45),
    .I0(x8_y50),
    .I1(x7_y45),
    .I2(1'b0),
    .I3(x8_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100111000000)
) lut_11_45 (
    .O(x11_y45),
    .I0(x9_y48),
    .I1(x8_y49),
    .I2(1'b0),
    .I3(x8_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011011100010)
) lut_12_45 (
    .O(x12_y45),
    .I0(x9_y46),
    .I1(x10_y44),
    .I2(x10_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000110111000)
) lut_13_45 (
    .O(x13_y45),
    .I0(x10_y47),
    .I1(x10_y43),
    .I2(1'b0),
    .I3(x10_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101011100101)
) lut_14_45 (
    .O(x14_y45),
    .I0(x12_y44),
    .I1(x11_y42),
    .I2(x12_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001110100011)
) lut_15_45 (
    .O(x15_y45),
    .I0(x12_y50),
    .I1(x13_y47),
    .I2(x13_y43),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111000110111)
) lut_16_45 (
    .O(x16_y45),
    .I0(x14_y48),
    .I1(x13_y49),
    .I2(1'b0),
    .I3(x14_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011100110011)
) lut_17_45 (
    .O(x17_y45),
    .I0(x15_y46),
    .I1(x15_y44),
    .I2(x14_y45),
    .I3(x14_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110001110001)
) lut_18_45 (
    .O(x18_y45),
    .I0(x16_y44),
    .I1(x16_y41),
    .I2(x16_y41),
    .I3(x15_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100111111011)
) lut_19_45 (
    .O(x19_y45),
    .I0(x16_y42),
    .I1(1'b0),
    .I2(x16_y50),
    .I3(x16_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101011001100)
) lut_20_45 (
    .O(x20_y45),
    .I0(x18_y40),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x18_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101111001010)
) lut_21_45 (
    .O(x21_y45),
    .I0(x19_y48),
    .I1(x18_y50),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010110100000)
) lut_22_45 (
    .O(x22_y45),
    .I0(x19_y48),
    .I1(x19_y41),
    .I2(1'b0),
    .I3(x19_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011011001111)
) lut_23_45 (
    .O(x23_y45),
    .I0(x20_y47),
    .I1(x20_y50),
    .I2(x20_y47),
    .I3(x20_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111010000100)
) lut_24_45 (
    .O(x24_y45),
    .I0(x22_y41),
    .I1(1'b0),
    .I2(x22_y49),
    .I3(x22_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000011101010)
) lut_25_45 (
    .O(x25_y45),
    .I0(x22_y42),
    .I1(x22_y40),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001011011010)
) lut_26_45 (
    .O(x26_y45),
    .I0(1'b0),
    .I1(x23_y42),
    .I2(1'b0),
    .I3(x24_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110010000110)
) lut_27_45 (
    .O(x27_y45),
    .I0(x25_y45),
    .I1(x25_y46),
    .I2(1'b0),
    .I3(x24_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100101001000)
) lut_28_45 (
    .O(x28_y45),
    .I0(1'b0),
    .I1(x26_y40),
    .I2(1'b0),
    .I3(x25_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101011101110)
) lut_29_45 (
    .O(x29_y45),
    .I0(x27_y46),
    .I1(1'b0),
    .I2(x27_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111101110101)
) lut_30_45 (
    .O(x30_y45),
    .I0(x28_y41),
    .I1(x28_y48),
    .I2(x28_y42),
    .I3(x27_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101011100011)
) lut_31_45 (
    .O(x31_y45),
    .I0(x29_y46),
    .I1(1'b0),
    .I2(x29_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110011111000)
) lut_32_45 (
    .O(x32_y45),
    .I0(x30_y47),
    .I1(1'b0),
    .I2(x30_y42),
    .I3(x29_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000010110011)
) lut_33_45 (
    .O(x33_y45),
    .I0(x30_y43),
    .I1(x31_y47),
    .I2(x31_y46),
    .I3(x30_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111001100010)
) lut_34_45 (
    .O(x34_y45),
    .I0(x32_y49),
    .I1(x32_y44),
    .I2(x31_y48),
    .I3(x32_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010111001010)
) lut_35_45 (
    .O(x35_y45),
    .I0(x33_y40),
    .I1(x32_y50),
    .I2(x33_y50),
    .I3(x33_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011110001100)
) lut_36_45 (
    .O(x36_y45),
    .I0(x34_y48),
    .I1(x34_y44),
    .I2(1'b0),
    .I3(x33_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110111100101)
) lut_37_45 (
    .O(x37_y45),
    .I0(x35_y50),
    .I1(x34_y40),
    .I2(x35_y40),
    .I3(x35_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101000101010)
) lut_38_45 (
    .O(x38_y45),
    .I0(x36_y47),
    .I1(x35_y43),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101000001111)
) lut_39_45 (
    .O(x39_y45),
    .I0(x37_y42),
    .I1(1'b0),
    .I2(x36_y46),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011100101110)
) lut_40_45 (
    .O(x40_y45),
    .I0(1'b0),
    .I1(x37_y48),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110101111010)
) lut_41_45 (
    .O(x41_y45),
    .I0(x38_y41),
    .I1(x38_y40),
    .I2(x39_y43),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101100011010)
) lut_42_45 (
    .O(x42_y45),
    .I0(x39_y49),
    .I1(x39_y42),
    .I2(x39_y49),
    .I3(x39_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000010001101)
) lut_43_45 (
    .O(x43_y45),
    .I0(x41_y45),
    .I1(1'b0),
    .I2(x40_y49),
    .I3(x41_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111010110110)
) lut_44_45 (
    .O(x44_y45),
    .I0(x41_y43),
    .I1(x41_y45),
    .I2(x41_y47),
    .I3(x42_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011100111111)
) lut_45_45 (
    .O(x45_y45),
    .I0(1'b0),
    .I1(x43_y47),
    .I2(x43_y45),
    .I3(x42_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000110011011)
) lut_46_45 (
    .O(x46_y45),
    .I0(x43_y46),
    .I1(x43_y45),
    .I2(x44_y41),
    .I3(x44_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100111100100)
) lut_47_45 (
    .O(x47_y45),
    .I0(x44_y48),
    .I1(x44_y42),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010111001110)
) lut_48_45 (
    .O(x48_y45),
    .I0(x46_y40),
    .I1(1'b0),
    .I2(x45_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111100111111)
) lut_49_45 (
    .O(x49_y45),
    .I0(x46_y46),
    .I1(x46_y43),
    .I2(1'b0),
    .I3(x47_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101001001001)
) lut_50_45 (
    .O(x50_y45),
    .I0(1'b0),
    .I1(x47_y47),
    .I2(x48_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010001111110)
) lut_51_45 (
    .O(x51_y45),
    .I0(x49_y47),
    .I1(x49_y41),
    .I2(x48_y43),
    .I3(x48_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000010110101)
) lut_52_45 (
    .O(x52_y45),
    .I0(1'b0),
    .I1(x50_y44),
    .I2(x50_y46),
    .I3(x49_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110110000001)
) lut_53_45 (
    .O(x53_y45),
    .I0(x51_y47),
    .I1(x50_y46),
    .I2(1'b0),
    .I3(x51_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010011111100)
) lut_54_45 (
    .O(x54_y45),
    .I0(1'b0),
    .I1(x52_y44),
    .I2(x52_y49),
    .I3(x51_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000100000111)
) lut_55_45 (
    .O(x55_y45),
    .I0(1'b0),
    .I1(x52_y48),
    .I2(x52_y48),
    .I3(x53_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111000101001)
) lut_56_45 (
    .O(x56_y45),
    .I0(x54_y48),
    .I1(x54_y41),
    .I2(x53_y40),
    .I3(x54_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011000100001)
) lut_57_45 (
    .O(x57_y45),
    .I0(x55_y42),
    .I1(x54_y49),
    .I2(1'b0),
    .I3(x55_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111111010001)
) lut_58_45 (
    .O(x58_y45),
    .I0(x56_y42),
    .I1(x56_y41),
    .I2(1'b0),
    .I3(x55_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111110111100)
) lut_59_45 (
    .O(x59_y45),
    .I0(x56_y40),
    .I1(x56_y49),
    .I2(1'b0),
    .I3(x57_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111000101001)
) lut_60_45 (
    .O(x60_y45),
    .I0(x58_y43),
    .I1(x57_y41),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100101101101)
) lut_61_45 (
    .O(x61_y45),
    .I0(x59_y50),
    .I1(x59_y42),
    .I2(x59_y41),
    .I3(x58_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101110001010)
) lut_62_45 (
    .O(x62_y45),
    .I0(1'b0),
    .I1(x59_y41),
    .I2(x59_y47),
    .I3(x60_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111011100101)
) lut_0_46 (
    .O(x0_y46),
    .I0(in6),
    .I1(1'b0),
    .I2(in0),
    .I3(in7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001100011111)
) lut_1_46 (
    .O(x1_y46),
    .I0(in4),
    .I1(1'b0),
    .I2(in0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111110101011)
) lut_2_46 (
    .O(x2_y46),
    .I0(1'b0),
    .I1(in8),
    .I2(in0),
    .I3(in4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001100110010)
) lut_3_46 (
    .O(x3_y46),
    .I0(in8),
    .I1(x1_y43),
    .I2(in6),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110101111011)
) lut_4_46 (
    .O(x4_y46),
    .I0(x2_y50),
    .I1(x2_y50),
    .I2(x1_y51),
    .I3(x2_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011101101101)
) lut_5_46 (
    .O(x5_y46),
    .I0(x3_y42),
    .I1(1'b0),
    .I2(x2_y50),
    .I3(x3_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111111011111)
) lut_6_46 (
    .O(x6_y46),
    .I0(x3_y47),
    .I1(x3_y42),
    .I2(x3_y41),
    .I3(x4_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001101110011)
) lut_7_46 (
    .O(x7_y46),
    .I0(x5_y43),
    .I1(x4_y51),
    .I2(x5_y47),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000000100000)
) lut_8_46 (
    .O(x8_y46),
    .I0(x6_y51),
    .I1(x5_y47),
    .I2(x6_y48),
    .I3(x6_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100010000110)
) lut_9_46 (
    .O(x9_y46),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x6_y48),
    .I3(x6_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010100111000)
) lut_10_46 (
    .O(x10_y46),
    .I0(x8_y49),
    .I1(1'b0),
    .I2(x8_y50),
    .I3(x8_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111001101110)
) lut_11_46 (
    .O(x11_y46),
    .I0(x9_y48),
    .I1(x9_y46),
    .I2(x8_y41),
    .I3(x9_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111111100100)
) lut_12_46 (
    .O(x12_y46),
    .I0(x9_y50),
    .I1(x10_y49),
    .I2(1'b0),
    .I3(x10_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100000010111)
) lut_13_46 (
    .O(x13_y46),
    .I0(x10_y48),
    .I1(x10_y41),
    .I2(x11_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100110010001)
) lut_14_46 (
    .O(x14_y46),
    .I0(x12_y41),
    .I1(x11_y42),
    .I2(x11_y44),
    .I3(x11_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011111110100)
) lut_15_46 (
    .O(x15_y46),
    .I0(x13_y41),
    .I1(x12_y43),
    .I2(x13_y41),
    .I3(x12_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101100110110)
) lut_16_46 (
    .O(x16_y46),
    .I0(x13_y45),
    .I1(x14_y51),
    .I2(x13_y41),
    .I3(x13_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011010000111)
) lut_17_46 (
    .O(x17_y46),
    .I0(x14_y47),
    .I1(x15_y48),
    .I2(x14_y46),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110100101100)
) lut_18_46 (
    .O(x18_y46),
    .I0(x16_y47),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x15_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010110010010)
) lut_19_46 (
    .O(x19_y46),
    .I0(x17_y46),
    .I1(x16_y47),
    .I2(x17_y47),
    .I3(x16_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011000010101)
) lut_20_46 (
    .O(x20_y46),
    .I0(x18_y42),
    .I1(x17_y47),
    .I2(x17_y41),
    .I3(x18_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000001100001)
) lut_21_46 (
    .O(x21_y46),
    .I0(x18_y48),
    .I1(x18_y43),
    .I2(x19_y48),
    .I3(x18_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101100001100)
) lut_22_46 (
    .O(x22_y46),
    .I0(x19_y42),
    .I1(1'b0),
    .I2(x20_y47),
    .I3(x20_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101010011110)
) lut_23_46 (
    .O(x23_y46),
    .I0(x21_y45),
    .I1(1'b0),
    .I2(x21_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011100100011)
) lut_24_46 (
    .O(x24_y46),
    .I0(x22_y51),
    .I1(1'b0),
    .I2(x22_y50),
    .I3(x21_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000110000000)
) lut_25_46 (
    .O(x25_y46),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x22_y45),
    .I3(x22_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001100110001)
) lut_26_46 (
    .O(x26_y46),
    .I0(x23_y48),
    .I1(x23_y49),
    .I2(x24_y50),
    .I3(x23_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011001011101)
) lut_27_46 (
    .O(x27_y46),
    .I0(x24_y50),
    .I1(1'b0),
    .I2(x25_y41),
    .I3(x25_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010000100110)
) lut_28_46 (
    .O(x28_y46),
    .I0(x25_y48),
    .I1(x26_y43),
    .I2(x25_y45),
    .I3(x26_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110010110110)
) lut_29_46 (
    .O(x29_y46),
    .I0(x27_y46),
    .I1(x27_y48),
    .I2(x26_y41),
    .I3(x27_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011100101001)
) lut_30_46 (
    .O(x30_y46),
    .I0(x28_y44),
    .I1(x27_y47),
    .I2(x27_y42),
    .I3(x28_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100101110111)
) lut_31_46 (
    .O(x31_y46),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x28_y48),
    .I3(x29_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110010101001)
) lut_32_46 (
    .O(x32_y46),
    .I0(x29_y50),
    .I1(x29_y42),
    .I2(x29_y45),
    .I3(x29_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000010111111)
) lut_33_46 (
    .O(x33_y46),
    .I0(1'b0),
    .I1(x31_y43),
    .I2(1'b0),
    .I3(x31_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110111001111)
) lut_34_46 (
    .O(x34_y46),
    .I0(x31_y51),
    .I1(x31_y46),
    .I2(x31_y49),
    .I3(x31_y41)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001011100000)
) lut_35_46 (
    .O(x35_y46),
    .I0(x33_y51),
    .I1(x32_y50),
    .I2(x33_y50),
    .I3(x33_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000001000010)
) lut_36_46 (
    .O(x36_y46),
    .I0(x34_y43),
    .I1(1'b0),
    .I2(x34_y41),
    .I3(x34_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011001111001)
) lut_37_46 (
    .O(x37_y46),
    .I0(1'b0),
    .I1(x35_y50),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010111001010)
) lut_38_46 (
    .O(x38_y46),
    .I0(x35_y50),
    .I1(1'b0),
    .I2(x36_y46),
    .I3(x35_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101001011010)
) lut_39_46 (
    .O(x39_y46),
    .I0(x37_y43),
    .I1(x36_y41),
    .I2(x37_y47),
    .I3(x37_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011110001010)
) lut_40_46 (
    .O(x40_y46),
    .I0(x37_y48),
    .I1(1'b0),
    .I2(x38_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111000001000)
) lut_41_46 (
    .O(x41_y46),
    .I0(x39_y51),
    .I1(x38_y47),
    .I2(x39_y43),
    .I3(x39_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100001110010)
) lut_42_46 (
    .O(x42_y46),
    .I0(x39_y45),
    .I1(x40_y45),
    .I2(x40_y41),
    .I3(x39_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111010001100)
) lut_43_46 (
    .O(x43_y46),
    .I0(x40_y43),
    .I1(x40_y50),
    .I2(x41_y50),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001100010101)
) lut_44_46 (
    .O(x44_y46),
    .I0(1'b0),
    .I1(x41_y44),
    .I2(x42_y47),
    .I3(x42_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001100101010)
) lut_45_46 (
    .O(x45_y46),
    .I0(x43_y51),
    .I1(x43_y48),
    .I2(1'b0),
    .I3(x42_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101111111111)
) lut_46_46 (
    .O(x46_y46),
    .I0(1'b0),
    .I1(x44_y44),
    .I2(x43_y41),
    .I3(x43_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111001011010)
) lut_47_46 (
    .O(x47_y46),
    .I0(x44_y45),
    .I1(x45_y43),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111000101011)
) lut_48_46 (
    .O(x48_y46),
    .I0(x45_y47),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x46_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101110110100)
) lut_49_46 (
    .O(x49_y46),
    .I0(1'b0),
    .I1(x46_y43),
    .I2(x46_y50),
    .I3(x47_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110100101111)
) lut_50_46 (
    .O(x50_y46),
    .I0(1'b0),
    .I1(x48_y42),
    .I2(x47_y46),
    .I3(x47_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010010101100)
) lut_51_46 (
    .O(x51_y46),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x49_y50),
    .I3(x48_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110100101011)
) lut_52_46 (
    .O(x52_y46),
    .I0(x50_y44),
    .I1(x49_y41),
    .I2(x49_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100011011110)
) lut_53_46 (
    .O(x53_y46),
    .I0(1'b0),
    .I1(x50_y44),
    .I2(x50_y45),
    .I3(x51_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000110100010)
) lut_54_46 (
    .O(x54_y46),
    .I0(x51_y45),
    .I1(x51_y41),
    .I2(x51_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011010100000)
) lut_55_46 (
    .O(x55_y46),
    .I0(x52_y45),
    .I1(x52_y50),
    .I2(x52_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111001100001)
) lut_56_46 (
    .O(x56_y46),
    .I0(x53_y43),
    .I1(x54_y41),
    .I2(x53_y43),
    .I3(x53_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100001101010)
) lut_57_46 (
    .O(x57_y46),
    .I0(1'b0),
    .I1(x55_y43),
    .I2(1'b0),
    .I3(x54_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101010010110)
) lut_58_46 (
    .O(x58_y46),
    .I0(x55_y41),
    .I1(x55_y44),
    .I2(x56_y46),
    .I3(x56_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101101111011)
) lut_59_46 (
    .O(x59_y46),
    .I0(x56_y41),
    .I1(x57_y51),
    .I2(x57_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011011011010)
) lut_60_46 (
    .O(x60_y46),
    .I0(x58_y49),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x57_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001101111101)
) lut_61_46 (
    .O(x61_y46),
    .I0(x59_y48),
    .I1(x59_y49),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101100100011)
) lut_62_46 (
    .O(x62_y46),
    .I0(1'b0),
    .I1(x60_y46),
    .I2(x60_y44),
    .I3(x59_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111000011101)
) lut_0_47 (
    .O(x0_y47),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(in4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101001010110)
) lut_1_47 (
    .O(x1_y47),
    .I0(in1),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100110111101)
) lut_2_47 (
    .O(x2_y47),
    .I0(in1),
    .I1(in2),
    .I2(in0),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010101100010)
) lut_3_47 (
    .O(x3_y47),
    .I0(in6),
    .I1(x1_y49),
    .I2(x1_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011110000001)
) lut_4_47 (
    .O(x4_y47),
    .I0(x2_y50),
    .I1(x1_y49),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100000110010)
) lut_5_47 (
    .O(x5_y47),
    .I0(1'b0),
    .I1(x3_y46),
    .I2(x2_y50),
    .I3(x2_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110100111110)
) lut_6_47 (
    .O(x6_y47),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x4_y49),
    .I3(x3_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111100101101)
) lut_7_47 (
    .O(x7_y47),
    .I0(x5_y48),
    .I1(x4_y46),
    .I2(x5_y47),
    .I3(x4_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000000001011)
) lut_8_47 (
    .O(x8_y47),
    .I0(x5_y51),
    .I1(x6_y44),
    .I2(x5_y45),
    .I3(x5_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100001101110)
) lut_9_47 (
    .O(x9_y47),
    .I0(x7_y43),
    .I1(x7_y51),
    .I2(x5_y45),
    .I3(x5_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100111100011)
) lut_10_47 (
    .O(x10_y47),
    .I0(x8_y47),
    .I1(x8_y45),
    .I2(x8_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111110111010)
) lut_11_47 (
    .O(x11_y47),
    .I0(x8_y46),
    .I1(x9_y44),
    .I2(1'b0),
    .I3(x9_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111100010110)
) lut_12_47 (
    .O(x12_y47),
    .I0(1'b0),
    .I1(x9_y48),
    .I2(1'b0),
    .I3(x9_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111001101101)
) lut_13_47 (
    .O(x13_y47),
    .I0(x10_y47),
    .I1(x10_y44),
    .I2(x11_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000100010000)
) lut_14_47 (
    .O(x14_y47),
    .I0(x11_y47),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x11_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111011101110)
) lut_15_47 (
    .O(x15_y47),
    .I0(x13_y47),
    .I1(x12_y52),
    .I2(x13_y48),
    .I3(x12_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011100010110)
) lut_16_47 (
    .O(x16_y47),
    .I0(x13_y47),
    .I1(1'b0),
    .I2(x13_y52),
    .I3(x14_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111010001000)
) lut_17_47 (
    .O(x17_y47),
    .I0(x15_y47),
    .I1(x15_y42),
    .I2(x15_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100110111111)
) lut_18_47 (
    .O(x18_y47),
    .I0(x15_y52),
    .I1(x15_y46),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011001011111)
) lut_19_47 (
    .O(x19_y47),
    .I0(1'b0),
    .I1(x16_y48),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000110010111)
) lut_20_47 (
    .O(x20_y47),
    .I0(x17_y45),
    .I1(x18_y52),
    .I2(x18_y48),
    .I3(x17_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100000001101)
) lut_21_47 (
    .O(x21_y47),
    .I0(x18_y42),
    .I1(x18_y42),
    .I2(1'b0),
    .I3(x19_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001011110001)
) lut_22_47 (
    .O(x22_y47),
    .I0(1'b0),
    .I1(x19_y43),
    .I2(x19_y50),
    .I3(x20_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110110100010)
) lut_23_47 (
    .O(x23_y47),
    .I0(x20_y42),
    .I1(1'b0),
    .I2(x20_y51),
    .I3(x20_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001100011011)
) lut_24_47 (
    .O(x24_y47),
    .I0(x21_y49),
    .I1(x22_y44),
    .I2(x21_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000010101100)
) lut_25_47 (
    .O(x25_y47),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x23_y44),
    .I3(x23_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100110110001)
) lut_26_47 (
    .O(x26_y47),
    .I0(x23_y44),
    .I1(1'b0),
    .I2(x23_y46),
    .I3(x24_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110011011000)
) lut_27_47 (
    .O(x27_y47),
    .I0(x25_y42),
    .I1(x24_y48),
    .I2(x24_y49),
    .I3(x24_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011000111110)
) lut_28_47 (
    .O(x28_y47),
    .I0(x25_y43),
    .I1(x25_y45),
    .I2(x25_y48),
    .I3(x26_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111011111010)
) lut_29_47 (
    .O(x29_y47),
    .I0(1'b0),
    .I1(x26_y47),
    .I2(x27_y43),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000100010110)
) lut_30_47 (
    .O(x30_y47),
    .I0(x27_y51),
    .I1(x27_y45),
    .I2(x27_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101000010001)
) lut_31_47 (
    .O(x31_y47),
    .I0(x29_y47),
    .I1(x29_y51),
    .I2(x28_y50),
    .I3(x28_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101100100101)
) lut_32_47 (
    .O(x32_y47),
    .I0(x30_y46),
    .I1(1'b0),
    .I2(x30_y44),
    .I3(x29_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101011101011)
) lut_33_47 (
    .O(x33_y47),
    .I0(x30_y47),
    .I1(x30_y48),
    .I2(x31_y49),
    .I3(x30_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000101100011)
) lut_34_47 (
    .O(x34_y47),
    .I0(x31_y49),
    .I1(x32_y51),
    .I2(x32_y52),
    .I3(x31_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110010001001)
) lut_35_47 (
    .O(x35_y47),
    .I0(x33_y52),
    .I1(x33_y51),
    .I2(1'b0),
    .I3(x32_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001101101111)
) lut_36_47 (
    .O(x36_y47),
    .I0(x33_y46),
    .I1(x33_y51),
    .I2(x34_y45),
    .I3(x34_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111011111110)
) lut_37_47 (
    .O(x37_y47),
    .I0(1'b0),
    .I1(x35_y47),
    .I2(x34_y49),
    .I3(x35_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110101011001)
) lut_38_47 (
    .O(x38_y47),
    .I0(1'b0),
    .I1(x35_y45),
    .I2(1'b0),
    .I3(x35_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001010010111)
) lut_39_47 (
    .O(x39_y47),
    .I0(x36_y51),
    .I1(x36_y45),
    .I2(x36_y50),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111000010101)
) lut_40_47 (
    .O(x40_y47),
    .I0(1'b0),
    .I1(x37_y46),
    .I2(1'b0),
    .I3(x38_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011000110110)
) lut_41_47 (
    .O(x41_y47),
    .I0(x38_y44),
    .I1(1'b0),
    .I2(x39_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110001101100)
) lut_42_47 (
    .O(x42_y47),
    .I0(x40_y44),
    .I1(1'b0),
    .I2(x40_y44),
    .I3(x40_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111110110011)
) lut_43_47 (
    .O(x43_y47),
    .I0(x40_y52),
    .I1(x40_y48),
    .I2(x40_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110110100001)
) lut_44_47 (
    .O(x44_y47),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x42_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110101001101)
) lut_45_47 (
    .O(x45_y47),
    .I0(x43_y50),
    .I1(x42_y50),
    .I2(x43_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100100111110)
) lut_46_47 (
    .O(x46_y47),
    .I0(x44_y48),
    .I1(x44_y51),
    .I2(x44_y47),
    .I3(x44_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110100010000)
) lut_47_47 (
    .O(x47_y47),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x45_y48),
    .I3(x44_y42)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101000010101)
) lut_48_47 (
    .O(x48_y47),
    .I0(x45_y49),
    .I1(x46_y42),
    .I2(x46_y48),
    .I3(x46_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001011100001)
) lut_49_47 (
    .O(x49_y47),
    .I0(x46_y44),
    .I1(x46_y42),
    .I2(x46_y49),
    .I3(x47_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101011011100)
) lut_50_47 (
    .O(x50_y47),
    .I0(x47_y44),
    .I1(x48_y51),
    .I2(x48_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111011011010)
) lut_51_47 (
    .O(x51_y47),
    .I0(x48_y48),
    .I1(x48_y44),
    .I2(x48_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101101110000)
) lut_52_47 (
    .O(x52_y47),
    .I0(x49_y49),
    .I1(x49_y47),
    .I2(x49_y49),
    .I3(x50_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010001011011)
) lut_53_47 (
    .O(x53_y47),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x51_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000011000111)
) lut_54_47 (
    .O(x54_y47),
    .I0(1'b0),
    .I1(x51_y45),
    .I2(x52_y42),
    .I3(x51_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100010100100)
) lut_55_47 (
    .O(x55_y47),
    .I0(x52_y43),
    .I1(1'b0),
    .I2(x53_y51),
    .I3(x52_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010000011110)
) lut_56_47 (
    .O(x56_y47),
    .I0(1'b0),
    .I1(x54_y46),
    .I2(x53_y42),
    .I3(x54_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110000011000)
) lut_57_47 (
    .O(x57_y47),
    .I0(x54_y46),
    .I1(x54_y48),
    .I2(x55_y52),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011101100011)
) lut_58_47 (
    .O(x58_y47),
    .I0(x55_y42),
    .I1(x56_y50),
    .I2(x55_y46),
    .I3(x55_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100111000000)
) lut_59_47 (
    .O(x59_y47),
    .I0(x56_y42),
    .I1(1'b0),
    .I2(x56_y44),
    .I3(x56_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110101100111)
) lut_60_47 (
    .O(x60_y47),
    .I0(x58_y45),
    .I1(x58_y50),
    .I2(x58_y44),
    .I3(x58_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000101101101)
) lut_61_47 (
    .O(x61_y47),
    .I0(1'b0),
    .I1(x59_y52),
    .I2(x58_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111011001011)
) lut_62_47 (
    .O(x62_y47),
    .I0(x60_y49),
    .I1(x60_y51),
    .I2(x60_y50),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111111010110)
) lut_0_48 (
    .O(x0_y48),
    .I0(1'b0),
    .I1(1'b0),
    .I2(in4),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001011010101)
) lut_1_48 (
    .O(x1_y48),
    .I0(in8),
    .I1(in5),
    .I2(in0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100000110101)
) lut_2_48 (
    .O(x2_y48),
    .I0(in3),
    .I1(in4),
    .I2(in4),
    .I3(in4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010011000010)
) lut_3_48 (
    .O(x3_y48),
    .I0(1'b0),
    .I1(x1_y43),
    .I2(in5),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011100111010)
) lut_4_48 (
    .O(x4_y48),
    .I0(1'b0),
    .I1(x1_y47),
    .I2(x1_y52),
    .I3(x1_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111001001011)
) lut_5_48 (
    .O(x5_y48),
    .I0(x2_y52),
    .I1(x2_y51),
    .I2(x2_y45),
    .I3(x3_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001001011011)
) lut_6_48 (
    .O(x6_y48),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x4_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101011101110)
) lut_7_48 (
    .O(x7_y48),
    .I0(x4_y49),
    .I1(x5_y47),
    .I2(x4_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101111110101)
) lut_8_48 (
    .O(x8_y48),
    .I0(1'b0),
    .I1(x6_y51),
    .I2(x6_y52),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000001111010)
) lut_9_48 (
    .O(x9_y48),
    .I0(1'b0),
    .I1(x7_y48),
    .I2(x6_y52),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101011000011)
) lut_10_48 (
    .O(x10_y48),
    .I0(x7_y48),
    .I1(x7_y44),
    .I2(x8_y45),
    .I3(x8_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111011111010)
) lut_11_48 (
    .O(x11_y48),
    .I0(1'b0),
    .I1(x8_y44),
    .I2(x8_y45),
    .I3(x8_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010001100001)
) lut_12_48 (
    .O(x12_y48),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x9_y51),
    .I3(x10_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010000101100)
) lut_13_48 (
    .O(x13_y48),
    .I0(1'b0),
    .I1(x11_y45),
    .I2(x10_y48),
    .I3(x10_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010100001001)
) lut_14_48 (
    .O(x14_y48),
    .I0(1'b0),
    .I1(x12_y48),
    .I2(x11_y53),
    .I3(x11_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011101011011)
) lut_15_48 (
    .O(x15_y48),
    .I0(x13_y47),
    .I1(x13_y46),
    .I2(1'b0),
    .I3(x13_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100001000001)
) lut_16_48 (
    .O(x16_y48),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x13_y51),
    .I3(x13_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010101001101)
) lut_17_48 (
    .O(x17_y48),
    .I0(x14_y51),
    .I1(x15_y49),
    .I2(x14_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010001001001)
) lut_18_48 (
    .O(x18_y48),
    .I0(x15_y47),
    .I1(1'b0),
    .I2(x15_y50),
    .I3(x15_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110011100111)
) lut_19_48 (
    .O(x19_y48),
    .I0(x16_y45),
    .I1(x16_y53),
    .I2(x17_y45),
    .I3(x17_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111111100011)
) lut_20_48 (
    .O(x20_y48),
    .I0(1'b0),
    .I1(x18_y51),
    .I2(x18_y49),
    .I3(x18_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110000111111)
) lut_21_48 (
    .O(x21_y48),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x18_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101011010001)
) lut_22_48 (
    .O(x22_y48),
    .I0(x19_y53),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x19_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011011000010)
) lut_23_48 (
    .O(x23_y48),
    .I0(1'b0),
    .I1(x21_y50),
    .I2(x21_y53),
    .I3(x20_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110010010101)
) lut_24_48 (
    .O(x24_y48),
    .I0(x22_y44),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x22_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100011100110)
) lut_25_48 (
    .O(x25_y48),
    .I0(x22_y47),
    .I1(x22_y45),
    .I2(1'b0),
    .I3(x23_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010000000010)
) lut_26_48 (
    .O(x26_y48),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x23_y53),
    .I3(x23_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000010011011)
) lut_27_48 (
    .O(x27_y48),
    .I0(x25_y46),
    .I1(x25_y47),
    .I2(x24_y51),
    .I3(x25_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100000100110)
) lut_28_48 (
    .O(x28_y48),
    .I0(1'b0),
    .I1(x26_y47),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011011100100)
) lut_29_48 (
    .O(x29_y48),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x27_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000001000101)
) lut_30_48 (
    .O(x30_y48),
    .I0(1'b0),
    .I1(x27_y51),
    .I2(x27_y47),
    .I3(x27_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000011000001)
) lut_31_48 (
    .O(x31_y48),
    .I0(x28_y52),
    .I1(x29_y44),
    .I2(x29_y53),
    .I3(x28_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111010011011)
) lut_32_48 (
    .O(x32_y48),
    .I0(x29_y52),
    .I1(x30_y49),
    .I2(1'b0),
    .I3(x29_y43)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100110001010)
) lut_33_48 (
    .O(x33_y48),
    .I0(x31_y46),
    .I1(x30_y50),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111100010010)
) lut_34_48 (
    .O(x34_y48),
    .I0(1'b0),
    .I1(x31_y51),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111000001001)
) lut_35_48 (
    .O(x35_y48),
    .I0(x33_y47),
    .I1(x32_y46),
    .I2(x33_y43),
    .I3(x32_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101101111001)
) lut_36_48 (
    .O(x36_y48),
    .I0(x33_y52),
    .I1(1'b0),
    .I2(x34_y46),
    .I3(x34_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011100110011)
) lut_37_48 (
    .O(x37_y48),
    .I0(x35_y46),
    .I1(x34_y53),
    .I2(x35_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010001001111)
) lut_38_48 (
    .O(x38_y48),
    .I0(x36_y53),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x35_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001100000111)
) lut_39_48 (
    .O(x39_y48),
    .I0(1'b0),
    .I1(x36_y53),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110111011111)
) lut_40_48 (
    .O(x40_y48),
    .I0(x38_y52),
    .I1(x37_y51),
    .I2(x37_y43),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100111111110)
) lut_41_48 (
    .O(x41_y48),
    .I0(x39_y44),
    .I1(x38_y52),
    .I2(x38_y50),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110101100111)
) lut_42_48 (
    .O(x42_y48),
    .I0(x40_y47),
    .I1(1'b0),
    .I2(x40_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110110101111)
) lut_43_48 (
    .O(x43_y48),
    .I0(x41_y45),
    .I1(1'b0),
    .I2(x40_y48),
    .I3(x40_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111010010011)
) lut_44_48 (
    .O(x44_y48),
    .I0(x42_y47),
    .I1(x42_y44),
    .I2(1'b0),
    .I3(x41_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111101011011)
) lut_45_48 (
    .O(x45_y48),
    .I0(x42_y46),
    .I1(x42_y52),
    .I2(x42_y45),
    .I3(x42_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110110010000)
) lut_46_48 (
    .O(x46_y48),
    .I0(x44_y48),
    .I1(x44_y46),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011001110010)
) lut_47_48 (
    .O(x47_y48),
    .I0(x44_y45),
    .I1(x44_y43),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110110010000)
) lut_48_48 (
    .O(x48_y48),
    .I0(x45_y45),
    .I1(x46_y44),
    .I2(x46_y44),
    .I3(x45_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101110011000)
) lut_49_48 (
    .O(x49_y48),
    .I0(x47_y48),
    .I1(x46_y47),
    .I2(x47_y53),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001111100010)
) lut_50_48 (
    .O(x50_y48),
    .I0(x47_y44),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101111011000)
) lut_51_48 (
    .O(x51_y48),
    .I0(x49_y53),
    .I1(x48_y47),
    .I2(x49_y50),
    .I3(x48_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000100100000)
) lut_52_48 (
    .O(x52_y48),
    .I0(x49_y51),
    .I1(x50_y43),
    .I2(x49_y52),
    .I3(x50_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000101100110)
) lut_53_48 (
    .O(x53_y48),
    .I0(x50_y45),
    .I1(x51_y52),
    .I2(x51_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101001000110)
) lut_54_48 (
    .O(x54_y48),
    .I0(x51_y46),
    .I1(x52_y52),
    .I2(x52_y47),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100111100001)
) lut_55_48 (
    .O(x55_y48),
    .I0(x52_y43),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x53_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110110111100)
) lut_56_48 (
    .O(x56_y48),
    .I0(x53_y46),
    .I1(x53_y53),
    .I2(1'b0),
    .I3(x53_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011010010110)
) lut_57_48 (
    .O(x57_y48),
    .I0(x54_y43),
    .I1(x54_y46),
    .I2(x55_y47),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100010111011)
) lut_58_48 (
    .O(x58_y48),
    .I0(x56_y47),
    .I1(1'b0),
    .I2(x55_y48),
    .I3(x56_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010010000111)
) lut_59_48 (
    .O(x59_y48),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x57_y51),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111011010101)
) lut_60_48 (
    .O(x60_y48),
    .I0(x58_y46),
    .I1(x58_y53),
    .I2(1'b0),
    .I3(x58_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101110000010)
) lut_61_48 (
    .O(x61_y48),
    .I0(x58_y53),
    .I1(x59_y46),
    .I2(x59_y46),
    .I3(x58_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011111011101)
) lut_62_48 (
    .O(x62_y48),
    .I0(1'b0),
    .I1(x60_y45),
    .I2(x59_y51),
    .I3(x59_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111110111011)
) lut_0_49 (
    .O(x0_y49),
    .I0(1'b0),
    .I1(in0),
    .I2(in6),
    .I3(in3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111100001111)
) lut_1_49 (
    .O(x1_y49),
    .I0(1'b0),
    .I1(in0),
    .I2(1'b0),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000011000000)
) lut_2_49 (
    .O(x2_y49),
    .I0(in4),
    .I1(in2),
    .I2(in1),
    .I3(in5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100111111011)
) lut_3_49 (
    .O(x3_y49),
    .I0(x1_y50),
    .I1(x1_y54),
    .I2(in3),
    .I3(in6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100010110011)
) lut_4_49 (
    .O(x4_y49),
    .I0(x2_y50),
    .I1(1'b0),
    .I2(x1_y50),
    .I3(x2_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001110110010)
) lut_5_49 (
    .O(x5_y49),
    .I0(x3_y48),
    .I1(x3_y45),
    .I2(x3_y52),
    .I3(x3_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100010101010)
) lut_6_49 (
    .O(x6_y49),
    .I0(x3_y48),
    .I1(x3_y47),
    .I2(x4_y50),
    .I3(x4_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111000100111)
) lut_7_49 (
    .O(x7_y49),
    .I0(x5_y54),
    .I1(x4_y47),
    .I2(1'b0),
    .I3(x5_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101010110011)
) lut_8_49 (
    .O(x8_y49),
    .I0(x6_y51),
    .I1(x5_y47),
    .I2(x5_y52),
    .I3(x6_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001110011010)
) lut_9_49 (
    .O(x9_y49),
    .I0(1'b0),
    .I1(x6_y54),
    .I2(x5_y52),
    .I3(x6_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011110001001)
) lut_10_49 (
    .O(x10_y49),
    .I0(x8_y49),
    .I1(x7_y50),
    .I2(x7_y44),
    .I3(x8_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001010001001)
) lut_11_49 (
    .O(x11_y49),
    .I0(x8_y52),
    .I1(x9_y54),
    .I2(x8_y54),
    .I3(x9_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101011000010)
) lut_12_49 (
    .O(x12_y49),
    .I0(x10_y51),
    .I1(1'b0),
    .I2(x10_y54),
    .I3(x10_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111010101001)
) lut_13_49 (
    .O(x13_y49),
    .I0(x10_y53),
    .I1(x10_y52),
    .I2(x11_y47),
    .I3(x10_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111100001011)
) lut_14_49 (
    .O(x14_y49),
    .I0(x12_y48),
    .I1(x11_y49),
    .I2(x12_y50),
    .I3(x11_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100110010111)
) lut_15_49 (
    .O(x15_y49),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x12_y49),
    .I3(x13_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001111001001)
) lut_16_49 (
    .O(x16_y49),
    .I0(x14_y50),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x13_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001001000010)
) lut_17_49 (
    .O(x17_y49),
    .I0(x15_y45),
    .I1(x15_y44),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000011000110)
) lut_18_49 (
    .O(x18_y49),
    .I0(1'b0),
    .I1(x15_y48),
    .I2(x16_y48),
    .I3(x15_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000011100010)
) lut_19_49 (
    .O(x19_y49),
    .I0(1'b0),
    .I1(x16_y44),
    .I2(x17_y53),
    .I3(x16_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101010000110)
) lut_20_49 (
    .O(x20_y49),
    .I0(x18_y49),
    .I1(x18_y46),
    .I2(1'b0),
    .I3(x18_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011100001000)
) lut_21_49 (
    .O(x21_y49),
    .I0(1'b0),
    .I1(x19_y49),
    .I2(1'b0),
    .I3(x19_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001111011010)
) lut_22_49 (
    .O(x22_y49),
    .I0(1'b0),
    .I1(x19_y49),
    .I2(x19_y48),
    .I3(x20_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010111010111)
) lut_23_49 (
    .O(x23_y49),
    .I0(x21_y45),
    .I1(x20_y53),
    .I2(x20_y51),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100100011101)
) lut_24_49 (
    .O(x24_y49),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x21_y54),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111010010010)
) lut_25_49 (
    .O(x25_y49),
    .I0(x22_y49),
    .I1(x22_y44),
    .I2(x23_y45),
    .I3(x23_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101101011111)
) lut_26_49 (
    .O(x26_y49),
    .I0(x24_y44),
    .I1(x24_y49),
    .I2(x24_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101010010111)
) lut_27_49 (
    .O(x27_y49),
    .I0(x25_y48),
    .I1(x24_y50),
    .I2(x25_y46),
    .I3(x24_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001011100111)
) lut_28_49 (
    .O(x28_y49),
    .I0(x26_y47),
    .I1(x26_y44),
    .I2(x25_y54),
    .I3(x26_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111100110010)
) lut_29_49 (
    .O(x29_y49),
    .I0(1'b0),
    .I1(x27_y54),
    .I2(x26_y45),
    .I3(x27_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111000010001)
) lut_30_49 (
    .O(x30_y49),
    .I0(x28_y49),
    .I1(x27_y47),
    .I2(x27_y52),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010101111100)
) lut_31_49 (
    .O(x31_y49),
    .I0(x29_y46),
    .I1(x29_y52),
    .I2(x28_y52),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110101010011)
) lut_32_49 (
    .O(x32_y49),
    .I0(x29_y51),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x29_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101000010010)
) lut_33_49 (
    .O(x33_y49),
    .I0(x31_y48),
    .I1(x31_y53),
    .I2(x31_y51),
    .I3(x31_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000000010100)
) lut_34_49 (
    .O(x34_y49),
    .I0(x32_y52),
    .I1(x31_y45),
    .I2(x31_y52),
    .I3(x31_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110011111001)
) lut_35_49 (
    .O(x35_y49),
    .I0(x32_y51),
    .I1(x33_y47),
    .I2(x32_y45),
    .I3(x33_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011001011000)
) lut_36_49 (
    .O(x36_y49),
    .I0(x34_y46),
    .I1(x34_y44),
    .I2(x34_y47),
    .I3(x33_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011111001111)
) lut_37_49 (
    .O(x37_y49),
    .I0(x35_y47),
    .I1(x35_y48),
    .I2(x34_y45),
    .I3(x35_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111100001100)
) lut_38_49 (
    .O(x38_y49),
    .I0(x36_y52),
    .I1(x35_y46),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100001110101)
) lut_39_49 (
    .O(x39_y49),
    .I0(x37_y50),
    .I1(1'b0),
    .I2(x37_y45),
    .I3(x37_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010101110101)
) lut_40_49 (
    .O(x40_y49),
    .I0(x38_y50),
    .I1(x38_y50),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100101100001)
) lut_41_49 (
    .O(x41_y49),
    .I0(x38_y53),
    .I1(x38_y49),
    .I2(x38_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001011101101)
) lut_42_49 (
    .O(x42_y49),
    .I0(x40_y48),
    .I1(x39_y52),
    .I2(x40_y49),
    .I3(x40_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101011110000)
) lut_43_49 (
    .O(x43_y49),
    .I0(x40_y48),
    .I1(x40_y54),
    .I2(x40_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111001100011)
) lut_44_49 (
    .O(x44_y49),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x41_y51),
    .I3(x42_y44)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100111010000)
) lut_45_49 (
    .O(x45_y49),
    .I0(1'b0),
    .I1(x42_y44),
    .I2(x43_y46),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111100001001)
) lut_46_49 (
    .O(x46_y49),
    .I0(x44_y52),
    .I1(x43_y49),
    .I2(x43_y46),
    .I3(x44_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111111010111)
) lut_47_49 (
    .O(x47_y49),
    .I0(x45_y50),
    .I1(x44_y45),
    .I2(x44_y53),
    .I3(x44_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001110001101)
) lut_48_49 (
    .O(x48_y49),
    .I0(x45_y49),
    .I1(x45_y51),
    .I2(x45_y54),
    .I3(x46_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100001110000)
) lut_49_49 (
    .O(x49_y49),
    .I0(x46_y50),
    .I1(x47_y52),
    .I2(x46_y48),
    .I3(x47_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001100101110)
) lut_50_49 (
    .O(x50_y49),
    .I0(x48_y45),
    .I1(x47_y47),
    .I2(x47_y50),
    .I3(x47_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010000011011)
) lut_51_49 (
    .O(x51_y49),
    .I0(x48_y48),
    .I1(x48_y53),
    .I2(x49_y47),
    .I3(x48_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001001010110)
) lut_52_49 (
    .O(x52_y49),
    .I0(x50_y44),
    .I1(x50_y54),
    .I2(1'b0),
    .I3(x49_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101001100011)
) lut_53_49 (
    .O(x53_y49),
    .I0(x51_y50),
    .I1(x51_y53),
    .I2(x50_y52),
    .I3(x50_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011001110000)
) lut_54_49 (
    .O(x54_y49),
    .I0(x52_y44),
    .I1(x52_y48),
    .I2(x51_y49),
    .I3(x52_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101011000001)
) lut_55_49 (
    .O(x55_y49),
    .I0(x53_y50),
    .I1(x53_y47),
    .I2(x53_y52),
    .I3(x52_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000111110011)
) lut_56_49 (
    .O(x56_y49),
    .I0(1'b0),
    .I1(x53_y45),
    .I2(x53_y47),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010010000010)
) lut_57_49 (
    .O(x57_y49),
    .I0(x55_y53),
    .I1(x54_y51),
    .I2(x55_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101110011101)
) lut_58_49 (
    .O(x58_y49),
    .I0(x55_y48),
    .I1(1'b0),
    .I2(x55_y52),
    .I3(x55_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101000000100)
) lut_59_49 (
    .O(x59_y49),
    .I0(x57_y46),
    .I1(x57_y45),
    .I2(x57_y54),
    .I3(x56_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100110010011)
) lut_60_49 (
    .O(x60_y49),
    .I0(x58_y54),
    .I1(x57_y48),
    .I2(1'b0),
    .I3(x57_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011011110101)
) lut_61_49 (
    .O(x61_y49),
    .I0(x58_y53),
    .I1(x59_y45),
    .I2(x59_y53),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000011000010)
) lut_62_49 (
    .O(x62_y49),
    .I0(x59_y47),
    .I1(x60_y46),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010110001110)
) lut_0_50 (
    .O(x0_y50),
    .I0(in6),
    .I1(in0),
    .I2(in9),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110100100110)
) lut_1_50 (
    .O(x1_y50),
    .I0(1'b0),
    .I1(1'b0),
    .I2(in5),
    .I3(in5)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110110111101)
) lut_2_50 (
    .O(x2_y50),
    .I0(in3),
    .I1(in4),
    .I2(in1),
    .I3(in9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011110000100)
) lut_3_50 (
    .O(x3_y50),
    .I0(1'b0),
    .I1(in0),
    .I2(in5),
    .I3(x1_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000010001111)
) lut_4_50 (
    .O(x4_y50),
    .I0(x2_y54),
    .I1(x2_y50),
    .I2(x2_y55),
    .I3(x2_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100001011110)
) lut_5_50 (
    .O(x5_y50),
    .I0(x2_y55),
    .I1(x3_y47),
    .I2(x3_y50),
    .I3(x2_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001001111000)
) lut_6_50 (
    .O(x6_y50),
    .I0(1'b0),
    .I1(x4_y46),
    .I2(x3_y45),
    .I3(x3_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110111111110)
) lut_7_50 (
    .O(x7_y50),
    .I0(1'b0),
    .I1(x4_y52),
    .I2(1'b0),
    .I3(x4_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100111111001)
) lut_8_50 (
    .O(x8_y50),
    .I0(1'b0),
    .I1(x6_y50),
    .I2(x5_y47),
    .I3(x5_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000010001110)
) lut_9_50 (
    .O(x9_y50),
    .I0(x7_y45),
    .I1(x6_y54),
    .I2(x5_y47),
    .I3(x5_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001101010000)
) lut_10_50 (
    .O(x10_y50),
    .I0(x8_y52),
    .I1(x7_y53),
    .I2(x7_y52),
    .I3(x7_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011001011100)
) lut_11_50 (
    .O(x11_y50),
    .I0(1'b0),
    .I1(x9_y55),
    .I2(x9_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001001011100)
) lut_12_50 (
    .O(x12_y50),
    .I0(1'b0),
    .I1(x10_y54),
    .I2(x10_y50),
    .I3(x9_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101100100110)
) lut_13_50 (
    .O(x13_y50),
    .I0(x10_y51),
    .I1(x10_y51),
    .I2(x10_y45),
    .I3(x10_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110010100100)
) lut_14_50 (
    .O(x14_y50),
    .I0(1'b0),
    .I1(x12_y50),
    .I2(x12_y48),
    .I3(x11_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010010110011)
) lut_15_50 (
    .O(x15_y50),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x13_y50),
    .I3(x13_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000000010010)
) lut_16_50 (
    .O(x16_y50),
    .I0(x14_y51),
    .I1(x13_y50),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101010100101)
) lut_17_50 (
    .O(x17_y50),
    .I0(x14_y55),
    .I1(x14_y52),
    .I2(x14_y47),
    .I3(x14_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100110100001)
) lut_18_50 (
    .O(x18_y50),
    .I0(x16_y54),
    .I1(x16_y48),
    .I2(x16_y53),
    .I3(x15_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010101101011)
) lut_19_50 (
    .O(x19_y50),
    .I0(x17_y55),
    .I1(1'b0),
    .I2(x16_y53),
    .I3(x17_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010000010011)
) lut_20_50 (
    .O(x20_y50),
    .I0(x17_y52),
    .I1(x17_y50),
    .I2(x17_y54),
    .I3(x17_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000100111100)
) lut_21_50 (
    .O(x21_y50),
    .I0(x19_y48),
    .I1(x18_y48),
    .I2(x19_y45),
    .I3(x18_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011010110001)
) lut_22_50 (
    .O(x22_y50),
    .I0(1'b0),
    .I1(x20_y53),
    .I2(x20_y53),
    .I3(x20_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010011011010)
) lut_23_50 (
    .O(x23_y50),
    .I0(x21_y45),
    .I1(x20_y51),
    .I2(1'b0),
    .I3(x20_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101111001101)
) lut_24_50 (
    .O(x24_y50),
    .I0(x22_y45),
    .I1(1'b0),
    .I2(x22_y50),
    .I3(x22_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100110101110)
) lut_25_50 (
    .O(x25_y50),
    .I0(x23_y47),
    .I1(1'b0),
    .I2(x23_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101110001101)
) lut_26_50 (
    .O(x26_y50),
    .I0(x24_y52),
    .I1(1'b0),
    .I2(x24_y48),
    .I3(x24_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010011011111)
) lut_27_50 (
    .O(x27_y50),
    .I0(x24_y53),
    .I1(x24_y48),
    .I2(x25_y46),
    .I3(x24_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001001111101)
) lut_28_50 (
    .O(x28_y50),
    .I0(1'b0),
    .I1(x26_y49),
    .I2(x25_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101011101010)
) lut_29_50 (
    .O(x29_y50),
    .I0(x26_y49),
    .I1(x26_y53),
    .I2(x26_y50),
    .I3(x27_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110101000010)
) lut_30_50 (
    .O(x30_y50),
    .I0(1'b0),
    .I1(x27_y47),
    .I2(1'b0),
    .I3(x27_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111100001111)
) lut_31_50 (
    .O(x31_y50),
    .I0(x29_y48),
    .I1(x28_y51),
    .I2(x28_y55),
    .I3(x28_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111011101001)
) lut_32_50 (
    .O(x32_y50),
    .I0(x30_y47),
    .I1(x29_y50),
    .I2(x30_y46),
    .I3(x30_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011010000111)
) lut_33_50 (
    .O(x33_y50),
    .I0(x31_y49),
    .I1(x31_y45),
    .I2(1'b0),
    .I3(x30_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110100111010)
) lut_34_50 (
    .O(x34_y50),
    .I0(x31_y53),
    .I1(x31_y50),
    .I2(x31_y50),
    .I3(x31_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010010100111)
) lut_35_50 (
    .O(x35_y50),
    .I0(x32_y45),
    .I1(x33_y52),
    .I2(x33_y52),
    .I3(x33_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100010000110)
) lut_36_50 (
    .O(x36_y50),
    .I0(1'b0),
    .I1(x33_y45),
    .I2(x34_y48),
    .I3(x34_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010011010010)
) lut_37_50 (
    .O(x37_y50),
    .I0(x34_y45),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x35_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100011111110)
) lut_38_50 (
    .O(x38_y50),
    .I0(x35_y48),
    .I1(1'b0),
    .I2(x35_y47),
    .I3(x35_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101100110001)
) lut_39_50 (
    .O(x39_y50),
    .I0(x37_y55),
    .I1(x37_y46),
    .I2(x36_y54),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010111100101)
) lut_40_50 (
    .O(x40_y50),
    .I0(1'b0),
    .I1(x37_y50),
    .I2(x38_y47),
    .I3(x37_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000101000101)
) lut_41_50 (
    .O(x41_y50),
    .I0(x39_y54),
    .I1(x38_y50),
    .I2(x39_y51),
    .I3(x39_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111010001110)
) lut_42_50 (
    .O(x42_y50),
    .I0(x40_y45),
    .I1(1'b0),
    .I2(x39_y55),
    .I3(x39_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111010100000)
) lut_43_50 (
    .O(x43_y50),
    .I0(x41_y48),
    .I1(x40_y52),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101101100010)
) lut_44_50 (
    .O(x44_y50),
    .I0(x42_y55),
    .I1(1'b0),
    .I2(x41_y50),
    .I3(x41_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111010010101)
) lut_45_50 (
    .O(x45_y50),
    .I0(x42_y48),
    .I1(x43_y52),
    .I2(x42_y54),
    .I3(x42_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000011101101)
) lut_46_50 (
    .O(x46_y50),
    .I0(x44_y52),
    .I1(x43_y46),
    .I2(x43_y47),
    .I3(x43_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011000101100)
) lut_47_50 (
    .O(x47_y50),
    .I0(x45_y45),
    .I1(x45_y50),
    .I2(x44_y46),
    .I3(x44_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000010001001)
) lut_48_50 (
    .O(x48_y50),
    .I0(x45_y46),
    .I1(1'b0),
    .I2(x46_y52),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001011111010)
) lut_49_50 (
    .O(x49_y50),
    .I0(x47_y51),
    .I1(x47_y51),
    .I2(1'b0),
    .I3(x46_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001011010010)
) lut_50_50 (
    .O(x50_y50),
    .I0(x47_y47),
    .I1(x48_y54),
    .I2(x47_y50),
    .I3(x47_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000110101010)
) lut_51_50 (
    .O(x51_y50),
    .I0(x49_y47),
    .I1(x48_y45),
    .I2(x48_y45),
    .I3(x49_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011111111101)
) lut_52_50 (
    .O(x52_y50),
    .I0(x50_y55),
    .I1(x50_y52),
    .I2(x49_y53),
    .I3(x50_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111101101011)
) lut_53_50 (
    .O(x53_y50),
    .I0(x51_y55),
    .I1(x50_y54),
    .I2(x50_y46),
    .I3(x51_y45)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011101110000)
) lut_54_50 (
    .O(x54_y50),
    .I0(x52_y46),
    .I1(x52_y52),
    .I2(x51_y49),
    .I3(x52_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010101000000)
) lut_55_50 (
    .O(x55_y50),
    .I0(x53_y47),
    .I1(x52_y50),
    .I2(x52_y47),
    .I3(x53_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111001011101)
) lut_56_50 (
    .O(x56_y50),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x54_y45),
    .I3(x53_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100011000111)
) lut_57_50 (
    .O(x57_y50),
    .I0(x54_y52),
    .I1(1'b0),
    .I2(x55_y54),
    .I3(x54_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011101000110)
) lut_58_50 (
    .O(x58_y50),
    .I0(1'b0),
    .I1(x55_y51),
    .I2(x55_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001011010101)
) lut_59_50 (
    .O(x59_y50),
    .I0(x57_y48),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110111100001)
) lut_60_50 (
    .O(x60_y50),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x58_y48),
    .I3(x58_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111000101100)
) lut_61_50 (
    .O(x61_y50),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x59_y53),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001110111010)
) lut_62_50 (
    .O(x62_y50),
    .I0(x59_y54),
    .I1(x59_y47),
    .I2(x60_y52),
    .I3(x59_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100011000000)
) lut_0_51 (
    .O(x0_y51),
    .I0(in7),
    .I1(in4),
    .I2(in2),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110110100101)
) lut_1_51 (
    .O(x1_y51),
    .I0(in6),
    .I1(1'b0),
    .I2(in1),
    .I3(in6)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011111000011)
) lut_2_51 (
    .O(x2_y51),
    .I0(in5),
    .I1(1'b0),
    .I2(in8),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000111111011)
) lut_3_51 (
    .O(x3_y51),
    .I0(x1_y49),
    .I1(x1_y51),
    .I2(in0),
    .I3(x1_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111110010110)
) lut_4_51 (
    .O(x4_y51),
    .I0(x2_y52),
    .I1(x1_y51),
    .I2(1'b0),
    .I3(x1_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110110100110)
) lut_5_51 (
    .O(x5_y51),
    .I0(x3_y47),
    .I1(x2_y47),
    .I2(1'b0),
    .I3(x3_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101001100110)
) lut_6_51 (
    .O(x6_y51),
    .I0(x4_y46),
    .I1(x4_y46),
    .I2(x4_y52),
    .I3(x4_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100110001000)
) lut_7_51 (
    .O(x7_y51),
    .I0(x4_y46),
    .I1(x4_y48),
    .I2(x5_y53),
    .I3(x4_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101001011001)
) lut_8_51 (
    .O(x8_y51),
    .I0(x5_y53),
    .I1(x6_y49),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100011100010)
) lut_9_51 (
    .O(x9_y51),
    .I0(x6_y47),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100111000100)
) lut_10_51 (
    .O(x10_y51),
    .I0(1'b0),
    .I1(x8_y47),
    .I2(x8_y49),
    .I3(x8_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111011111111)
) lut_11_51 (
    .O(x11_y51),
    .I0(x8_y54),
    .I1(x9_y56),
    .I2(1'b0),
    .I3(x8_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000110111010)
) lut_12_51 (
    .O(x12_y51),
    .I0(x9_y55),
    .I1(x9_y48),
    .I2(x10_y50),
    .I3(x9_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000001100111)
) lut_13_51 (
    .O(x13_y51),
    .I0(x11_y56),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x10_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110001011001)
) lut_14_51 (
    .O(x14_y51),
    .I0(x12_y55),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x12_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001000100000)
) lut_15_51 (
    .O(x15_y51),
    .I0(x12_y49),
    .I1(1'b0),
    .I2(x12_y54),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000011001010)
) lut_16_51 (
    .O(x16_y51),
    .I0(x14_y55),
    .I1(x13_y47),
    .I2(x13_y48),
    .I3(x13_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111000001100)
) lut_17_51 (
    .O(x17_y51),
    .I0(1'b0),
    .I1(x15_y47),
    .I2(x14_y50),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100000011011)
) lut_18_51 (
    .O(x18_y51),
    .I0(x15_y52),
    .I1(x15_y46),
    .I2(x15_y56),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111010111100)
) lut_19_51 (
    .O(x19_y51),
    .I0(x16_y46),
    .I1(1'b0),
    .I2(x16_y55),
    .I3(x17_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001101100101)
) lut_20_51 (
    .O(x20_y51),
    .I0(x17_y51),
    .I1(1'b0),
    .I2(x18_y47),
    .I3(x18_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100110000110)
) lut_21_51 (
    .O(x21_y51),
    .I0(x19_y47),
    .I1(x19_y51),
    .I2(1'b0),
    .I3(x18_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001010101010)
) lut_22_51 (
    .O(x22_y51),
    .I0(x19_y54),
    .I1(x20_y53),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011110100111)
) lut_23_51 (
    .O(x23_y51),
    .I0(1'b0),
    .I1(x21_y55),
    .I2(x20_y55),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101011010100)
) lut_24_51 (
    .O(x24_y51),
    .I0(x21_y48),
    .I1(x22_y54),
    .I2(x22_y55),
    .I3(x21_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101100000010)
) lut_25_51 (
    .O(x25_y51),
    .I0(x23_y56),
    .I1(x22_y52),
    .I2(x22_y49),
    .I3(x22_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110100000010)
) lut_26_51 (
    .O(x26_y51),
    .I0(x23_y56),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x24_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111010111110)
) lut_27_51 (
    .O(x27_y51),
    .I0(x25_y46),
    .I1(x25_y56),
    .I2(x25_y52),
    .I3(x25_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001001101011)
) lut_28_51 (
    .O(x28_y51),
    .I0(1'b0),
    .I1(x25_y48),
    .I2(x25_y47),
    .I3(x25_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000010001101)
) lut_29_51 (
    .O(x29_y51),
    .I0(x26_y46),
    .I1(x27_y53),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101100001011)
) lut_30_51 (
    .O(x30_y51),
    .I0(x28_y52),
    .I1(1'b0),
    .I2(x27_y53),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010110011001)
) lut_31_51 (
    .O(x31_y51),
    .I0(x29_y52),
    .I1(x29_y47),
    .I2(1'b0),
    .I3(x29_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100000110101)
) lut_32_51 (
    .O(x32_y51),
    .I0(x29_y51),
    .I1(x29_y47),
    .I2(1'b0),
    .I3(x29_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100000100111)
) lut_33_51 (
    .O(x33_y51),
    .I0(x31_y48),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x31_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011000110000)
) lut_34_51 (
    .O(x34_y51),
    .I0(x31_y52),
    .I1(x32_y47),
    .I2(x31_y50),
    .I3(x31_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111000010100)
) lut_35_51 (
    .O(x35_y51),
    .I0(x33_y50),
    .I1(x33_y56),
    .I2(x33_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111011000000)
) lut_36_51 (
    .O(x36_y51),
    .I0(x33_y54),
    .I1(x33_y50),
    .I2(1'b0),
    .I3(x33_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110010110011)
) lut_37_51 (
    .O(x37_y51),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x35_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010001111110)
) lut_38_51 (
    .O(x38_y51),
    .I0(x36_y56),
    .I1(1'b0),
    .I2(x36_y55),
    .I3(x35_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011011011011)
) lut_39_51 (
    .O(x39_y51),
    .I0(1'b0),
    .I1(x36_y49),
    .I2(x37_y56),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000101101000)
) lut_40_51 (
    .O(x40_y51),
    .I0(x37_y51),
    .I1(x38_y47),
    .I2(x37_y48),
    .I3(x37_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000011101100)
) lut_41_51 (
    .O(x41_y51),
    .I0(1'b0),
    .I1(x38_y48),
    .I2(x38_y56),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110010110100)
) lut_42_51 (
    .O(x42_y51),
    .I0(x40_y49),
    .I1(x39_y56),
    .I2(1'b0),
    .I3(x39_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111010011101)
) lut_43_51 (
    .O(x43_y51),
    .I0(x41_y53),
    .I1(1'b0),
    .I2(x41_y50),
    .I3(x41_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010000111101)
) lut_44_51 (
    .O(x44_y51),
    .I0(x42_y52),
    .I1(1'b0),
    .I2(x41_y56),
    .I3(x41_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100111101010)
) lut_45_51 (
    .O(x45_y51),
    .I0(1'b0),
    .I1(x42_y48),
    .I2(1'b0),
    .I3(x43_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000000001010)
) lut_46_51 (
    .O(x46_y51),
    .I0(1'b0),
    .I1(x44_y48),
    .I2(x43_y55),
    .I3(x44_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001010010100)
) lut_47_51 (
    .O(x47_y51),
    .I0(x44_y55),
    .I1(1'b0),
    .I2(x44_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100111100000)
) lut_48_51 (
    .O(x48_y51),
    .I0(1'b0),
    .I1(x45_y55),
    .I2(x46_y55),
    .I3(x46_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001110111111)
) lut_49_51 (
    .O(x49_y51),
    .I0(x46_y54),
    .I1(x46_y54),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010111010110)
) lut_50_51 (
    .O(x50_y51),
    .I0(x47_y47),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010010111001)
) lut_51_51 (
    .O(x51_y51),
    .I0(1'b0),
    .I1(x49_y48),
    .I2(1'b0),
    .I3(x49_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100001001010)
) lut_52_51 (
    .O(x52_y51),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x49_y55),
    .I3(x49_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011111110010)
) lut_53_51 (
    .O(x53_y51),
    .I0(1'b0),
    .I1(x51_y47),
    .I2(x50_y54),
    .I3(x50_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000010100111)
) lut_54_51 (
    .O(x54_y51),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x52_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001101010101)
) lut_55_51 (
    .O(x55_y51),
    .I0(x52_y48),
    .I1(x52_y52),
    .I2(x52_y49),
    .I3(x53_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110001011011)
) lut_56_51 (
    .O(x56_y51),
    .I0(x53_y49),
    .I1(x53_y54),
    .I2(x53_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000000111110)
) lut_57_51 (
    .O(x57_y51),
    .I0(x54_y55),
    .I1(x55_y52),
    .I2(1'b0),
    .I3(x54_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010101010111)
) lut_58_51 (
    .O(x58_y51),
    .I0(x56_y53),
    .I1(1'b0),
    .I2(x55_y48),
    .I3(x56_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110101111001)
) lut_59_51 (
    .O(x59_y51),
    .I0(x57_y54),
    .I1(1'b0),
    .I2(x57_y54),
    .I3(x56_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000001010111)
) lut_60_51 (
    .O(x60_y51),
    .I0(x57_y47),
    .I1(x58_y51),
    .I2(x57_y50),
    .I3(x58_y46)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010111110000)
) lut_61_51 (
    .O(x61_y51),
    .I0(x58_y47),
    .I1(1'b0),
    .I2(x58_y47),
    .I3(x58_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101100101000)
) lut_62_51 (
    .O(x62_y51),
    .I0(x59_y56),
    .I1(1'b0),
    .I2(x60_y52),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110101110011)
) lut_0_52 (
    .O(x0_y52),
    .I0(in3),
    .I1(in4),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100100001101)
) lut_1_52 (
    .O(x1_y52),
    .I0(in0),
    .I1(1'b0),
    .I2(in7),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100000000001)
) lut_2_52 (
    .O(x2_y52),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(in3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101000001001)
) lut_3_52 (
    .O(x3_y52),
    .I0(1'b0),
    .I1(x1_y47),
    .I2(in0),
    .I3(x1_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111101110111)
) lut_4_52 (
    .O(x4_y52),
    .I0(x2_y57),
    .I1(x1_y47),
    .I2(x2_y52),
    .I3(x2_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000101100101)
) lut_5_52 (
    .O(x5_y52),
    .I0(x3_y48),
    .I1(x3_y52),
    .I2(x2_y56),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011111111010)
) lut_6_52 (
    .O(x6_y52),
    .I0(x3_y51),
    .I1(x3_y52),
    .I2(x3_y57),
    .I3(x4_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011001111101)
) lut_7_52 (
    .O(x7_y52),
    .I0(x4_y47),
    .I1(1'b0),
    .I2(x4_y49),
    .I3(x4_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011001011111)
) lut_8_52 (
    .O(x8_y52),
    .I0(x6_y47),
    .I1(x5_y56),
    .I2(x5_y56),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011010011001)
) lut_9_52 (
    .O(x9_y52),
    .I0(x7_y49),
    .I1(x7_y48),
    .I2(x5_y56),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100100000001)
) lut_10_52 (
    .O(x10_y52),
    .I0(x7_y53),
    .I1(x8_y50),
    .I2(x7_y47),
    .I3(x7_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110110010100)
) lut_11_52 (
    .O(x11_y52),
    .I0(x9_y53),
    .I1(x9_y48),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110110100100)
) lut_12_52 (
    .O(x12_y52),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x9_y57),
    .I3(x9_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111010101111)
) lut_13_52 (
    .O(x13_y52),
    .I0(x11_y56),
    .I1(x10_y50),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001001001010)
) lut_14_52 (
    .O(x14_y52),
    .I0(1'b0),
    .I1(x11_y50),
    .I2(x12_y55),
    .I3(x11_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111010010010)
) lut_15_52 (
    .O(x15_y52),
    .I0(x12_y54),
    .I1(x13_y54),
    .I2(x13_y49),
    .I3(x13_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100001001110)
) lut_16_52 (
    .O(x16_y52),
    .I0(x14_y57),
    .I1(x13_y53),
    .I2(1'b0),
    .I3(x14_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000101000000)
) lut_17_52 (
    .O(x17_y52),
    .I0(1'b0),
    .I1(x14_y53),
    .I2(x14_y51),
    .I3(x14_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101000000010)
) lut_18_52 (
    .O(x18_y52),
    .I0(1'b0),
    .I1(x16_y50),
    .I2(x16_y55),
    .I3(x15_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010000111001)
) lut_19_52 (
    .O(x19_y52),
    .I0(x17_y54),
    .I1(x16_y53),
    .I2(x16_y51),
    .I3(x16_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110111100000)
) lut_20_52 (
    .O(x20_y52),
    .I0(x18_y47),
    .I1(x18_y51),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110001011100)
) lut_21_52 (
    .O(x21_y52),
    .I0(x19_y55),
    .I1(x18_y48),
    .I2(x18_y50),
    .I3(x18_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010011110000)
) lut_22_52 (
    .O(x22_y52),
    .I0(1'b0),
    .I1(x19_y52),
    .I2(x19_y55),
    .I3(x19_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011000000101)
) lut_23_52 (
    .O(x23_y52),
    .I0(x21_y47),
    .I1(x20_y47),
    .I2(x21_y55),
    .I3(x20_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010011111101)
) lut_24_52 (
    .O(x24_y52),
    .I0(x22_y54),
    .I1(x21_y50),
    .I2(x22_y57),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100000110001)
) lut_25_52 (
    .O(x25_y52),
    .I0(x23_y54),
    .I1(1'b0),
    .I2(x22_y55),
    .I3(x22_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011111001000)
) lut_26_52 (
    .O(x26_y52),
    .I0(x24_y56),
    .I1(x24_y56),
    .I2(x23_y53),
    .I3(x24_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100100001100)
) lut_27_52 (
    .O(x27_y52),
    .I0(x25_y48),
    .I1(x24_y50),
    .I2(1'b0),
    .I3(x25_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001010001110)
) lut_28_52 (
    .O(x28_y52),
    .I0(x25_y54),
    .I1(x25_y56),
    .I2(x25_y55),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010100110100)
) lut_29_52 (
    .O(x29_y52),
    .I0(x26_y47),
    .I1(x26_y50),
    .I2(x26_y54),
    .I3(x27_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001111001011)
) lut_30_52 (
    .O(x30_y52),
    .I0(x28_y50),
    .I1(x28_y54),
    .I2(1'b0),
    .I3(x27_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001101110110)
) lut_31_52 (
    .O(x31_y52),
    .I0(x28_y52),
    .I1(x28_y54),
    .I2(1'b0),
    .I3(x28_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011001001101)
) lut_32_52 (
    .O(x32_y52),
    .I0(1'b0),
    .I1(x29_y49),
    .I2(x30_y51),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110000111010)
) lut_33_52 (
    .O(x33_y52),
    .I0(1'b0),
    .I1(x31_y48),
    .I2(x30_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100001000001)
) lut_34_52 (
    .O(x34_y52),
    .I0(x31_y57),
    .I1(x32_y55),
    .I2(x32_y47),
    .I3(x32_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001010101101)
) lut_35_52 (
    .O(x35_y52),
    .I0(x32_y53),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000100111111)
) lut_36_52 (
    .O(x36_y52),
    .I0(1'b0),
    .I1(x33_y56),
    .I2(x33_y56),
    .I3(x34_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100100001100)
) lut_37_52 (
    .O(x37_y52),
    .I0(1'b0),
    .I1(x34_y50),
    .I2(x35_y52),
    .I3(x35_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011001100010)
) lut_38_52 (
    .O(x38_y52),
    .I0(x35_y56),
    .I1(1'b0),
    .I2(x35_y56),
    .I3(x36_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111000110000)
) lut_39_52 (
    .O(x39_y52),
    .I0(x36_y52),
    .I1(x37_y53),
    .I2(x37_y56),
    .I3(x36_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000000100100)
) lut_40_52 (
    .O(x40_y52),
    .I0(x37_y54),
    .I1(x37_y48),
    .I2(x38_y57),
    .I3(x37_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001110100000)
) lut_41_52 (
    .O(x41_y52),
    .I0(x39_y50),
    .I1(x39_y57),
    .I2(x38_y55),
    .I3(x39_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010101111111)
) lut_42_52 (
    .O(x42_y52),
    .I0(x39_y47),
    .I1(x40_y53),
    .I2(x39_y54),
    .I3(x39_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101000011100)
) lut_43_52 (
    .O(x43_y52),
    .I0(x40_y56),
    .I1(x41_y54),
    .I2(x40_y54),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111011100101)
) lut_44_52 (
    .O(x44_y52),
    .I0(x42_y48),
    .I1(x41_y54),
    .I2(x41_y51),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111110110001)
) lut_45_52 (
    .O(x45_y52),
    .I0(x42_y56),
    .I1(x43_y52),
    .I2(x43_y49),
    .I3(x42_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000000111001)
) lut_46_52 (
    .O(x46_y52),
    .I0(x44_y55),
    .I1(1'b0),
    .I2(x44_y50),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000110101011)
) lut_47_52 (
    .O(x47_y52),
    .I0(x45_y48),
    .I1(1'b0),
    .I2(x45_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011000100100)
) lut_48_52 (
    .O(x48_y52),
    .I0(x46_y51),
    .I1(1'b0),
    .I2(x45_y55),
    .I3(x46_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111011101000)
) lut_49_52 (
    .O(x49_y52),
    .I0(1'b0),
    .I1(x46_y47),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011111101111)
) lut_50_52 (
    .O(x50_y52),
    .I0(x48_y55),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x47_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000111111100)
) lut_51_52 (
    .O(x51_y52),
    .I0(x49_y57),
    .I1(x48_y52),
    .I2(x48_y53),
    .I3(x49_y47)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110111110101)
) lut_52_52 (
    .O(x52_y52),
    .I0(1'b0),
    .I1(x50_y55),
    .I2(x50_y51),
    .I3(x49_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000110111000)
) lut_53_52 (
    .O(x53_y52),
    .I0(1'b0),
    .I1(x50_y51),
    .I2(x50_y49),
    .I3(x50_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110010000101)
) lut_54_52 (
    .O(x54_y52),
    .I0(x52_y50),
    .I1(x52_y57),
    .I2(x52_y49),
    .I3(x52_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010001000011)
) lut_55_52 (
    .O(x55_y52),
    .I0(x52_y50),
    .I1(x52_y57),
    .I2(1'b0),
    .I3(x53_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101111001110)
) lut_56_52 (
    .O(x56_y52),
    .I0(1'b0),
    .I1(x54_y49),
    .I2(x53_y57),
    .I3(x53_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001110101100)
) lut_57_52 (
    .O(x57_y52),
    .I0(1'b0),
    .I1(x55_y54),
    .I2(x55_y49),
    .I3(x55_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101000001011)
) lut_58_52 (
    .O(x58_y52),
    .I0(1'b0),
    .I1(x55_y48),
    .I2(x55_y54),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001111110011)
) lut_59_52 (
    .O(x59_y52),
    .I0(x57_y52),
    .I1(1'b0),
    .I2(x57_y55),
    .I3(x56_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011110101110)
) lut_60_52 (
    .O(x60_y52),
    .I0(x57_y51),
    .I1(x58_y48),
    .I2(x58_y49),
    .I3(x58_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010111110001)
) lut_61_52 (
    .O(x61_y52),
    .I0(1'b0),
    .I1(x58_y49),
    .I2(x59_y56),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110010000011)
) lut_62_52 (
    .O(x62_y52),
    .I0(x59_y48),
    .I1(x59_y54),
    .I2(x60_y56),
    .I3(x59_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001101001101)
) lut_0_53 (
    .O(x0_y53),
    .I0(1'b0),
    .I1(in0),
    .I2(in0),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110011101100)
) lut_1_53 (
    .O(x1_y53),
    .I0(in4),
    .I1(in2),
    .I2(in6),
    .I3(in3)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101110010101)
) lut_2_53 (
    .O(x2_y53),
    .I0(in6),
    .I1(1'b0),
    .I2(in8),
    .I3(in9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010110111111)
) lut_3_53 (
    .O(x3_y53),
    .I0(in0),
    .I1(in0),
    .I2(in1),
    .I3(x1_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101111100111)
) lut_4_53 (
    .O(x4_y53),
    .I0(x1_y57),
    .I1(x1_y53),
    .I2(x1_y51),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011100111000)
) lut_5_53 (
    .O(x5_y53),
    .I0(x2_y53),
    .I1(x2_y54),
    .I2(x2_y56),
    .I3(x2_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011010000110)
) lut_6_53 (
    .O(x6_y53),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x3_y55),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101010100011)
) lut_7_53 (
    .O(x7_y53),
    .I0(x5_y48),
    .I1(1'b0),
    .I2(x4_y49),
    .I3(x4_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110000000100)
) lut_8_53 (
    .O(x8_y53),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x6_y49),
    .I3(x6_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101100010010)
) lut_9_53 (
    .O(x9_y53),
    .I0(x6_y53),
    .I1(1'b0),
    .I2(x6_y49),
    .I3(x6_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010101000101)
) lut_10_53 (
    .O(x10_y53),
    .I0(1'b0),
    .I1(x8_y58),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011101010000)
) lut_11_53 (
    .O(x11_y53),
    .I0(x8_y51),
    .I1(x9_y53),
    .I2(x8_y58),
    .I3(x8_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110101101100)
) lut_12_53 (
    .O(x12_y53),
    .I0(1'b0),
    .I1(x10_y52),
    .I2(x9_y51),
    .I3(x10_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011100001001)
) lut_13_53 (
    .O(x13_y53),
    .I0(x11_y58),
    .I1(1'b0),
    .I2(x10_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010100011001)
) lut_14_53 (
    .O(x14_y53),
    .I0(x11_y55),
    .I1(x11_y58),
    .I2(x11_y52),
    .I3(x11_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100111000001)
) lut_15_53 (
    .O(x15_y53),
    .I0(1'b0),
    .I1(x13_y49),
    .I2(1'b0),
    .I3(x12_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111110010100)
) lut_16_53 (
    .O(x16_y53),
    .I0(x14_y58),
    .I1(x13_y49),
    .I2(x14_y56),
    .I3(x13_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001011010110)
) lut_17_53 (
    .O(x17_y53),
    .I0(x15_y56),
    .I1(x15_y57),
    .I2(1'b0),
    .I3(x15_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001111001011)
) lut_18_53 (
    .O(x18_y53),
    .I0(x16_y57),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x15_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111100001011)
) lut_19_53 (
    .O(x19_y53),
    .I0(x17_y53),
    .I1(x16_y51),
    .I2(x16_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000101001110)
) lut_20_53 (
    .O(x20_y53),
    .I0(x18_y48),
    .I1(1'b0),
    .I2(x18_y49),
    .I3(x17_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011110100101)
) lut_21_53 (
    .O(x21_y53),
    .I0(1'b0),
    .I1(x19_y49),
    .I2(x18_y58),
    .I3(x19_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011000001100)
) lut_22_53 (
    .O(x22_y53),
    .I0(x19_y58),
    .I1(x20_y56),
    .I2(x19_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000010110110)
) lut_23_53 (
    .O(x23_y53),
    .I0(x21_y58),
    .I1(x21_y58),
    .I2(x20_y49),
    .I3(x20_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111100010110)
) lut_24_53 (
    .O(x24_y53),
    .I0(1'b0),
    .I1(x22_y48),
    .I2(x21_y57),
    .I3(x21_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010010100101)
) lut_25_53 (
    .O(x25_y53),
    .I0(x22_y53),
    .I1(x23_y48),
    .I2(x23_y53),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011101001010)
) lut_26_53 (
    .O(x26_y53),
    .I0(1'b0),
    .I1(x24_y57),
    .I2(x23_y50),
    .I3(x23_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110010000100)
) lut_27_53 (
    .O(x27_y53),
    .I0(x24_y54),
    .I1(x24_y54),
    .I2(x24_y49),
    .I3(x25_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011110000111)
) lut_28_53 (
    .O(x28_y53),
    .I0(1'b0),
    .I1(x26_y54),
    .I2(x25_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010001101001)
) lut_29_53 (
    .O(x29_y53),
    .I0(x26_y53),
    .I1(x27_y58),
    .I2(1'b0),
    .I3(x26_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101000101011)
) lut_30_53 (
    .O(x30_y53),
    .I0(x28_y54),
    .I1(x27_y58),
    .I2(x28_y48),
    .I3(x28_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110001110110)
) lut_31_53 (
    .O(x31_y53),
    .I0(x29_y51),
    .I1(x29_y57),
    .I2(1'b0),
    .I3(x28_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110111110010)
) lut_32_53 (
    .O(x32_y53),
    .I0(x29_y48),
    .I1(1'b0),
    .I2(x30_y56),
    .I3(x30_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111110010101)
) lut_33_53 (
    .O(x33_y53),
    .I0(x30_y58),
    .I1(x31_y48),
    .I2(x31_y48),
    .I3(x30_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000110101111)
) lut_34_53 (
    .O(x34_y53),
    .I0(x32_y57),
    .I1(1'b0),
    .I2(x32_y51),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100001101101)
) lut_35_53 (
    .O(x35_y53),
    .I0(x32_y58),
    .I1(x32_y52),
    .I2(x33_y51),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011010110010)
) lut_36_53 (
    .O(x36_y53),
    .I0(1'b0),
    .I1(x34_y50),
    .I2(x33_y50),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000010011101)
) lut_37_53 (
    .O(x37_y53),
    .I0(x35_y56),
    .I1(1'b0),
    .I2(x34_y49),
    .I3(x35_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001011100110)
) lut_38_53 (
    .O(x38_y53),
    .I0(x36_y51),
    .I1(x36_y56),
    .I2(1'b0),
    .I3(x36_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001110011011)
) lut_39_53 (
    .O(x39_y53),
    .I0(x37_y58),
    .I1(x36_y51),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011111001010)
) lut_40_53 (
    .O(x40_y53),
    .I0(x37_y49),
    .I1(x37_y50),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101101001101)
) lut_41_53 (
    .O(x41_y53),
    .I0(x39_y56),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x39_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111001111010)
) lut_42_53 (
    .O(x42_y53),
    .I0(1'b0),
    .I1(x40_y50),
    .I2(x40_y54),
    .I3(x40_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101011000001)
) lut_43_53 (
    .O(x43_y53),
    .I0(1'b0),
    .I1(x41_y51),
    .I2(x40_y51),
    .I3(x41_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111000111001)
) lut_44_53 (
    .O(x44_y53),
    .I0(x41_y50),
    .I1(x41_y54),
    .I2(1'b0),
    .I3(x42_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111011011101)
) lut_45_53 (
    .O(x45_y53),
    .I0(x42_y56),
    .I1(x43_y50),
    .I2(1'b0),
    .I3(x42_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000110101010)
) lut_46_53 (
    .O(x46_y53),
    .I0(x44_y48),
    .I1(x43_y57),
    .I2(x43_y53),
    .I3(x43_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000101101101)
) lut_47_53 (
    .O(x47_y53),
    .I0(x45_y50),
    .I1(x44_y48),
    .I2(x45_y54),
    .I3(x44_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101110010011)
) lut_48_53 (
    .O(x48_y53),
    .I0(x45_y49),
    .I1(x45_y57),
    .I2(x46_y55),
    .I3(x45_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011000100010)
) lut_49_53 (
    .O(x49_y53),
    .I0(x47_y52),
    .I1(x46_y58),
    .I2(1'b0),
    .I3(x47_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011111100111)
) lut_50_53 (
    .O(x50_y53),
    .I0(x48_y49),
    .I1(x48_y48),
    .I2(x48_y58),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000010000111)
) lut_51_53 (
    .O(x51_y53),
    .I0(x48_y55),
    .I1(x49_y50),
    .I2(x48_y48),
    .I3(x48_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011001111111)
) lut_52_53 (
    .O(x52_y53),
    .I0(x50_y54),
    .I1(x50_y55),
    .I2(x50_y57),
    .I3(x50_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011100011100)
) lut_53_53 (
    .O(x53_y53),
    .I0(1'b0),
    .I1(x50_y48),
    .I2(1'b0),
    .I3(x51_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101111010110)
) lut_54_53 (
    .O(x54_y53),
    .I0(1'b0),
    .I1(x52_y55),
    .I2(x51_y57),
    .I3(x52_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101011100001)
) lut_55_53 (
    .O(x55_y53),
    .I0(1'b0),
    .I1(x53_y54),
    .I2(x52_y49),
    .I3(x52_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101100001011)
) lut_56_53 (
    .O(x56_y53),
    .I0(x53_y54),
    .I1(x54_y51),
    .I2(1'b0),
    .I3(x53_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111111101001)
) lut_57_53 (
    .O(x57_y53),
    .I0(x55_y48),
    .I1(x55_y54),
    .I2(x55_y51),
    .I3(x55_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000011101101)
) lut_58_53 (
    .O(x58_y53),
    .I0(1'b0),
    .I1(x56_y49),
    .I2(x56_y57),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001111111100)
) lut_59_53 (
    .O(x59_y53),
    .I0(x56_y49),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x57_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100001110100)
) lut_60_53 (
    .O(x60_y53),
    .I0(x58_y50),
    .I1(x58_y52),
    .I2(x58_y52),
    .I3(x58_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111000010110)
) lut_61_53 (
    .O(x61_y53),
    .I0(x59_y54),
    .I1(x58_y58),
    .I2(x59_y52),
    .I3(x59_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111110000101)
) lut_62_53 (
    .O(x62_y53),
    .I0(x60_y50),
    .I1(1'b0),
    .I2(x60_y51),
    .I3(x59_y48)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101110011100)
) lut_0_54 (
    .O(x0_y54),
    .I0(in5),
    .I1(in4),
    .I2(in9),
    .I3(in9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100111011010)
) lut_1_54 (
    .O(x1_y54),
    .I0(in9),
    .I1(in8),
    .I2(in5),
    .I3(in4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111000100101)
) lut_2_54 (
    .O(x2_y54),
    .I0(1'b0),
    .I1(in4),
    .I2(1'b0),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000100010101)
) lut_3_54 (
    .O(x3_y54),
    .I0(1'b0),
    .I1(x1_y50),
    .I2(x1_y56),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101010011011)
) lut_4_54 (
    .O(x4_y54),
    .I0(1'b0),
    .I1(x1_y57),
    .I2(x2_y52),
    .I3(x2_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110111011001)
) lut_5_54 (
    .O(x5_y54),
    .I0(x3_y55),
    .I1(x2_y52),
    .I2(x3_y50),
    .I3(x2_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001011001100)
) lut_6_54 (
    .O(x6_y54),
    .I0(1'b0),
    .I1(x4_y58),
    .I2(x4_y50),
    .I3(x3_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000110010110)
) lut_7_54 (
    .O(x7_y54),
    .I0(x5_y50),
    .I1(x5_y51),
    .I2(x4_y51),
    .I3(x4_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001010110001)
) lut_8_54 (
    .O(x8_y54),
    .I0(x5_y51),
    .I1(x6_y57),
    .I2(1'b0),
    .I3(x6_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110100110010)
) lut_9_54 (
    .O(x9_y54),
    .I0(x7_y56),
    .I1(x7_y49),
    .I2(1'b0),
    .I3(x6_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011001110100)
) lut_10_54 (
    .O(x10_y54),
    .I0(x8_y57),
    .I1(1'b0),
    .I2(x7_y58),
    .I3(x7_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110100011000)
) lut_11_54 (
    .O(x11_y54),
    .I0(x9_y54),
    .I1(x8_y50),
    .I2(1'b0),
    .I3(x9_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010101001111)
) lut_12_54 (
    .O(x12_y54),
    .I0(x9_y50),
    .I1(x9_y51),
    .I2(1'b0),
    .I3(x9_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000000001100)
) lut_13_54 (
    .O(x13_y54),
    .I0(1'b0),
    .I1(x11_y54),
    .I2(x10_y53),
    .I3(x11_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101001010111)
) lut_14_54 (
    .O(x14_y54),
    .I0(x12_y49),
    .I1(x12_y52),
    .I2(x11_y58),
    .I3(x12_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011111101000)
) lut_15_54 (
    .O(x15_y54),
    .I0(x13_y49),
    .I1(x13_y56),
    .I2(x12_y51),
    .I3(x12_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010010011001)
) lut_16_54 (
    .O(x16_y54),
    .I0(x13_y53),
    .I1(x14_y55),
    .I2(1'b0),
    .I3(x14_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001101101110)
) lut_17_54 (
    .O(x17_y54),
    .I0(1'b0),
    .I1(x14_y49),
    .I2(x15_y53),
    .I3(x14_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010111110111)
) lut_18_54 (
    .O(x18_y54),
    .I0(x16_y53),
    .I1(x15_y52),
    .I2(x15_y56),
    .I3(x16_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111011101001)
) lut_19_54 (
    .O(x19_y54),
    .I0(x17_y59),
    .I1(1'b0),
    .I2(x17_y58),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001110011011)
) lut_20_54 (
    .O(x20_y54),
    .I0(x17_y55),
    .I1(1'b0),
    .I2(x18_y58),
    .I3(x17_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000001100001)
) lut_21_54 (
    .O(x21_y54),
    .I0(x19_y59),
    .I1(1'b0),
    .I2(x18_y59),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101010110101)
) lut_22_54 (
    .O(x22_y54),
    .I0(1'b0),
    .I1(x20_y50),
    .I2(x20_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001101011000)
) lut_23_54 (
    .O(x23_y54),
    .I0(1'b0),
    .I1(x20_y53),
    .I2(x21_y55),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111101100001)
) lut_24_54 (
    .O(x24_y54),
    .I0(1'b0),
    .I1(x21_y57),
    .I2(x22_y51),
    .I3(x22_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100111110100)
) lut_25_54 (
    .O(x25_y54),
    .I0(x23_y53),
    .I1(1'b0),
    .I2(x23_y56),
    .I3(x22_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101101011011)
) lut_26_54 (
    .O(x26_y54),
    .I0(x23_y52),
    .I1(x23_y53),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101101101010)
) lut_27_54 (
    .O(x27_y54),
    .I0(x24_y58),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x24_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000100010100)
) lut_28_54 (
    .O(x28_y54),
    .I0(x25_y55),
    .I1(x25_y58),
    .I2(x26_y59),
    .I3(x26_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100100001111)
) lut_29_54 (
    .O(x29_y54),
    .I0(x27_y55),
    .I1(x26_y51),
    .I2(x26_y53),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101000000100)
) lut_30_54 (
    .O(x30_y54),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x27_y49),
    .I3(x27_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110000010001)
) lut_31_54 (
    .O(x31_y54),
    .I0(x28_y51),
    .I1(x29_y52),
    .I2(x28_y54),
    .I3(x29_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100110101011)
) lut_32_54 (
    .O(x32_y54),
    .I0(x29_y55),
    .I1(x29_y56),
    .I2(x29_y51),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110110010001)
) lut_33_54 (
    .O(x33_y54),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x30_y52),
    .I3(x30_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100010111010)
) lut_34_54 (
    .O(x34_y54),
    .I0(x32_y56),
    .I1(x32_y53),
    .I2(x32_y58),
    .I3(x31_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101100101111)
) lut_35_54 (
    .O(x35_y54),
    .I0(1'b0),
    .I1(x32_y50),
    .I2(x33_y59),
    .I3(x32_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100111010111)
) lut_36_54 (
    .O(x36_y54),
    .I0(1'b0),
    .I1(x33_y57),
    .I2(x33_y49),
    .I3(x34_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100101111001)
) lut_37_54 (
    .O(x37_y54),
    .I0(x34_y51),
    .I1(x34_y55),
    .I2(x35_y51),
    .I3(x34_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110100010000)
) lut_38_54 (
    .O(x38_y54),
    .I0(1'b0),
    .I1(x35_y55),
    .I2(x35_y50),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111011100110)
) lut_39_54 (
    .O(x39_y54),
    .I0(1'b0),
    .I1(x36_y56),
    .I2(x37_y52),
    .I3(x37_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100001100110)
) lut_40_54 (
    .O(x40_y54),
    .I0(x38_y49),
    .I1(x37_y50),
    .I2(x38_y58),
    .I3(x38_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001001010101)
) lut_41_54 (
    .O(x41_y54),
    .I0(x39_y53),
    .I1(x38_y59),
    .I2(x38_y55),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111000010010)
) lut_42_54 (
    .O(x42_y54),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x39_y59),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011011110011)
) lut_43_54 (
    .O(x43_y54),
    .I0(1'b0),
    .I1(x40_y59),
    .I2(x40_y51),
    .I3(x41_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011100011101)
) lut_44_54 (
    .O(x44_y54),
    .I0(x41_y58),
    .I1(x42_y50),
    .I2(x41_y50),
    .I3(x42_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011001101010)
) lut_45_54 (
    .O(x45_y54),
    .I0(x42_y50),
    .I1(x43_y49),
    .I2(1'b0),
    .I3(x43_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100000011100)
) lut_46_54 (
    .O(x46_y54),
    .I0(1'b0),
    .I1(x43_y54),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101111000010)
) lut_47_54 (
    .O(x47_y54),
    .I0(x44_y58),
    .I1(x45_y59),
    .I2(x45_y59),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101101111110)
) lut_48_54 (
    .O(x48_y54),
    .I0(x46_y57),
    .I1(x46_y49),
    .I2(x45_y54),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011011000111)
) lut_49_54 (
    .O(x49_y54),
    .I0(x47_y55),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x46_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101100011110)
) lut_50_54 (
    .O(x50_y54),
    .I0(x47_y53),
    .I1(x47_y56),
    .I2(x48_y53),
    .I3(x48_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101110011111)
) lut_51_54 (
    .O(x51_y54),
    .I0(x49_y54),
    .I1(x49_y58),
    .I2(x48_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010111110011)
) lut_52_54 (
    .O(x52_y54),
    .I0(x49_y57),
    .I1(x50_y58),
    .I2(x49_y50),
    .I3(x49_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111010000100)
) lut_53_54 (
    .O(x53_y54),
    .I0(x50_y49),
    .I1(1'b0),
    .I2(x50_y49),
    .I3(x50_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000011100011)
) lut_54_54 (
    .O(x54_y54),
    .I0(x52_y51),
    .I1(x51_y59),
    .I2(x51_y56),
    .I3(x51_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001000001001)
) lut_55_54 (
    .O(x55_y54),
    .I0(x52_y50),
    .I1(x52_y59),
    .I2(x53_y55),
    .I3(x52_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010011010001)
) lut_56_54 (
    .O(x56_y54),
    .I0(x53_y55),
    .I1(x54_y53),
    .I2(x54_y59),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110001110100)
) lut_57_54 (
    .O(x57_y54),
    .I0(x55_y57),
    .I1(1'b0),
    .I2(x55_y59),
    .I3(x55_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110001010011)
) lut_58_54 (
    .O(x58_y54),
    .I0(x56_y56),
    .I1(x56_y51),
    .I2(x56_y56),
    .I3(x56_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100111111000)
) lut_59_54 (
    .O(x59_y54),
    .I0(x57_y56),
    .I1(x56_y51),
    .I2(x57_y53),
    .I3(x56_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010011110011)
) lut_60_54 (
    .O(x60_y54),
    .I0(x57_y51),
    .I1(x57_y56),
    .I2(x58_y55),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011010001111)
) lut_61_54 (
    .O(x61_y54),
    .I0(x59_y57),
    .I1(1'b0),
    .I2(x58_y54),
    .I3(x58_y49)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000100110100)
) lut_62_54 (
    .O(x62_y54),
    .I0(x60_y57),
    .I1(x60_y52),
    .I2(x60_y55),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011110011100)
) lut_0_55 (
    .O(x0_y55),
    .I0(in8),
    .I1(1'b0),
    .I2(in7),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001101110101)
) lut_1_55 (
    .O(x1_y55),
    .I0(1'b0),
    .I1(1'b0),
    .I2(in4),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010110011100)
) lut_2_55 (
    .O(x2_y55),
    .I0(in7),
    .I1(in8),
    .I2(in4),
    .I3(in9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111100001000)
) lut_3_55 (
    .O(x3_y55),
    .I0(x1_y59),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101011010101)
) lut_4_55 (
    .O(x4_y55),
    .I0(1'b0),
    .I1(x2_y53),
    .I2(x2_y60),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101000101010)
) lut_5_55 (
    .O(x5_y55),
    .I0(x3_y52),
    .I1(x3_y59),
    .I2(x2_y53),
    .I3(x2_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001111110001)
) lut_6_55 (
    .O(x6_y55),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x3_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010000110100)
) lut_7_55 (
    .O(x7_y55),
    .I0(x5_y56),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x4_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110110110110)
) lut_8_55 (
    .O(x8_y55),
    .I0(1'b0),
    .I1(x6_y50),
    .I2(x5_y59),
    .I3(x6_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110000110110)
) lut_9_55 (
    .O(x9_y55),
    .I0(x6_y58),
    .I1(x6_y50),
    .I2(x5_y59),
    .I3(x6_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000010010100)
) lut_10_55 (
    .O(x10_y55),
    .I0(x8_y50),
    .I1(x7_y60),
    .I2(x7_y50),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101001000000)
) lut_11_55 (
    .O(x11_y55),
    .I0(x8_y59),
    .I1(x9_y51),
    .I2(x8_y55),
    .I3(x8_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111100011101)
) lut_12_55 (
    .O(x12_y55),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x9_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101010001111)
) lut_13_55 (
    .O(x13_y55),
    .I0(x11_y50),
    .I1(x11_y52),
    .I2(x10_y53),
    .I3(x10_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101011111100)
) lut_14_55 (
    .O(x14_y55),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x12_y50),
    .I3(x12_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100011010001)
) lut_15_55 (
    .O(x15_y55),
    .I0(1'b0),
    .I1(x12_y54),
    .I2(x12_y52),
    .I3(x13_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001111011011)
) lut_16_55 (
    .O(x16_y55),
    .I0(x13_y53),
    .I1(x14_y54),
    .I2(x13_y50),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111000100001)
) lut_17_55 (
    .O(x17_y55),
    .I0(x14_y60),
    .I1(x15_y56),
    .I2(x14_y55),
    .I3(x15_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010111010010)
) lut_18_55 (
    .O(x18_y55),
    .I0(x15_y52),
    .I1(1'b0),
    .I2(x15_y50),
    .I3(x16_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011001001111)
) lut_19_55 (
    .O(x19_y55),
    .I0(1'b0),
    .I1(x16_y57),
    .I2(x17_y57),
    .I3(x17_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010111001100)
) lut_20_55 (
    .O(x20_y55),
    .I0(1'b0),
    .I1(x17_y51),
    .I2(1'b0),
    .I3(x17_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110110001111)
) lut_21_55 (
    .O(x21_y55),
    .I0(x19_y52),
    .I1(x18_y56),
    .I2(x19_y57),
    .I3(x18_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011011010011)
) lut_22_55 (
    .O(x22_y55),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101110001011)
) lut_23_55 (
    .O(x23_y55),
    .I0(x21_y50),
    .I1(x20_y51),
    .I2(x21_y56),
    .I3(x20_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000011011000)
) lut_24_55 (
    .O(x24_y55),
    .I0(x22_y54),
    .I1(x22_y51),
    .I2(x22_y54),
    .I3(x21_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000110010001)
) lut_25_55 (
    .O(x25_y55),
    .I0(x23_y60),
    .I1(1'b0),
    .I2(x22_y51),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000001100110)
) lut_26_55 (
    .O(x26_y55),
    .I0(x24_y58),
    .I1(1'b0),
    .I2(x24_y55),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011001011011)
) lut_27_55 (
    .O(x27_y55),
    .I0(x25_y57),
    .I1(x24_y57),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000101010101)
) lut_28_55 (
    .O(x28_y55),
    .I0(1'b0),
    .I1(x26_y50),
    .I2(x26_y51),
    .I3(x25_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100110011100)
) lut_29_55 (
    .O(x29_y55),
    .I0(x27_y57),
    .I1(x26_y50),
    .I2(x26_y55),
    .I3(x26_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110111011010)
) lut_30_55 (
    .O(x30_y55),
    .I0(x28_y60),
    .I1(x27_y59),
    .I2(x28_y52),
    .I3(x28_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111010010111)
) lut_31_55 (
    .O(x31_y55),
    .I0(x29_y56),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x29_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011110010111)
) lut_32_55 (
    .O(x32_y55),
    .I0(x29_y55),
    .I1(x30_y60),
    .I2(x30_y52),
    .I3(x29_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010010110001)
) lut_33_55 (
    .O(x33_y55),
    .I0(x31_y54),
    .I1(x31_y59),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101010001011)
) lut_34_55 (
    .O(x34_y55),
    .I0(x32_y52),
    .I1(x31_y59),
    .I2(x32_y60),
    .I3(x32_y50)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110011111010)
) lut_35_55 (
    .O(x35_y55),
    .I0(x33_y60),
    .I1(x32_y60),
    .I2(x33_y52),
    .I3(x32_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110100111011)
) lut_36_55 (
    .O(x36_y55),
    .I0(1'b0),
    .I1(x33_y57),
    .I2(x34_y51),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000100001110)
) lut_37_55 (
    .O(x37_y55),
    .I0(x35_y59),
    .I1(x35_y58),
    .I2(x34_y50),
    .I3(x35_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000011101001)
) lut_38_55 (
    .O(x38_y55),
    .I0(x36_y55),
    .I1(x36_y55),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000100010110)
) lut_39_55 (
    .O(x39_y55),
    .I0(x37_y57),
    .I1(x36_y52),
    .I2(x36_y54),
    .I3(x36_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101110010100)
) lut_40_55 (
    .O(x40_y55),
    .I0(x38_y54),
    .I1(x38_y54),
    .I2(x37_y51),
    .I3(x37_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100010111000)
) lut_41_55 (
    .O(x41_y55),
    .I0(1'b0),
    .I1(x38_y60),
    .I2(x38_y57),
    .I3(x38_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001101000110)
) lut_42_55 (
    .O(x42_y55),
    .I0(x40_y52),
    .I1(1'b0),
    .I2(x39_y56),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101101111110)
) lut_43_55 (
    .O(x43_y55),
    .I0(x41_y52),
    .I1(x41_y50),
    .I2(x40_y50),
    .I3(x41_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011110011100)
) lut_44_55 (
    .O(x44_y55),
    .I0(x42_y50),
    .I1(x42_y51),
    .I2(x41_y59),
    .I3(x42_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011111100010)
) lut_45_55 (
    .O(x45_y55),
    .I0(x43_y52),
    .I1(x43_y53),
    .I2(x43_y60),
    .I3(x42_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000101101000)
) lut_46_55 (
    .O(x46_y55),
    .I0(x44_y54),
    .I1(1'b0),
    .I2(x43_y54),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100101111001)
) lut_47_55 (
    .O(x47_y55),
    .I0(x45_y60),
    .I1(x45_y59),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011010000011)
) lut_48_55 (
    .O(x48_y55),
    .I0(x45_y50),
    .I1(1'b0),
    .I2(x46_y51),
    .I3(x46_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101010011000)
) lut_49_55 (
    .O(x49_y55),
    .I0(x47_y54),
    .I1(1'b0),
    .I2(x47_y60),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110111010011)
) lut_50_55 (
    .O(x50_y55),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x47_y58),
    .I3(x48_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101100010100)
) lut_51_55 (
    .O(x51_y55),
    .I0(x48_y53),
    .I1(1'b0),
    .I2(x49_y52),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000111101010)
) lut_52_55 (
    .O(x52_y55),
    .I0(x49_y60),
    .I1(x50_y52),
    .I2(1'b0),
    .I3(x49_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011000001010)
) lut_53_55 (
    .O(x53_y55),
    .I0(x50_y56),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x50_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110011011110)
) lut_54_55 (
    .O(x54_y55),
    .I0(x51_y54),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x51_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011110111100)
) lut_55_55 (
    .O(x55_y55),
    .I0(x52_y59),
    .I1(x53_y55),
    .I2(x52_y59),
    .I3(x53_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010000111100)
) lut_56_55 (
    .O(x56_y55),
    .I0(1'b0),
    .I1(x54_y60),
    .I2(x54_y54),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010100100010)
) lut_57_55 (
    .O(x57_y55),
    .I0(x55_y60),
    .I1(x55_y56),
    .I2(x54_y50),
    .I3(x54_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100110110100)
) lut_58_55 (
    .O(x58_y55),
    .I0(1'b0),
    .I1(x56_y53),
    .I2(x55_y58),
    .I3(x56_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001010101010)
) lut_59_55 (
    .O(x59_y55),
    .I0(x57_y53),
    .I1(x56_y57),
    .I2(x56_y56),
    .I3(x57_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110101000011)
) lut_60_55 (
    .O(x60_y55),
    .I0(x57_y57),
    .I1(x58_y56),
    .I2(x58_y52),
    .I3(x58_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101101100101)
) lut_61_55 (
    .O(x61_y55),
    .I0(x59_y57),
    .I1(1'b0),
    .I2(x58_y58),
    .I3(x58_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001010000010)
) lut_62_55 (
    .O(x62_y55),
    .I0(x59_y52),
    .I1(x60_y54),
    .I2(x60_y60),
    .I3(x59_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111100110110)
) lut_0_56 (
    .O(x0_y56),
    .I0(in0),
    .I1(in9),
    .I2(1'b0),
    .I3(in1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001010011111)
) lut_1_56 (
    .O(x1_y56),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(in9)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001101001100)
) lut_2_56 (
    .O(x2_y56),
    .I0(in8),
    .I1(in1),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111111110010)
) lut_3_56 (
    .O(x3_y56),
    .I0(x1_y60),
    .I1(x1_y52),
    .I2(in1),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001110100111)
) lut_4_56 (
    .O(x4_y56),
    .I0(x1_y59),
    .I1(x2_y53),
    .I2(x2_y60),
    .I3(x1_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010011011100)
) lut_5_56 (
    .O(x5_y56),
    .I0(x3_y58),
    .I1(x3_y61),
    .I2(x3_y58),
    .I3(x2_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001010111111)
) lut_6_56 (
    .O(x6_y56),
    .I0(1'b0),
    .I1(x3_y60),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101011000111)
) lut_7_56 (
    .O(x7_y56),
    .I0(x5_y60),
    .I1(x4_y58),
    .I2(x5_y60),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010000111000)
) lut_8_56 (
    .O(x8_y56),
    .I0(1'b0),
    .I1(x6_y57),
    .I2(x6_y57),
    .I3(x6_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110011000011)
) lut_9_56 (
    .O(x9_y56),
    .I0(x6_y55),
    .I1(1'b0),
    .I2(x6_y57),
    .I3(x6_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011111011010)
) lut_10_56 (
    .O(x10_y56),
    .I0(x7_y56),
    .I1(x8_y52),
    .I2(x7_y55),
    .I3(x8_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011010001010)
) lut_11_56 (
    .O(x11_y56),
    .I0(x9_y60),
    .I1(x8_y51),
    .I2(x8_y54),
    .I3(x9_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110100001111)
) lut_12_56 (
    .O(x12_y56),
    .I0(x9_y60),
    .I1(x10_y56),
    .I2(1'b0),
    .I3(x9_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000010111011)
) lut_13_56 (
    .O(x13_y56),
    .I0(x11_y60),
    .I1(x10_y57),
    .I2(x11_y61),
    .I3(x10_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000010111010)
) lut_14_56 (
    .O(x14_y56),
    .I0(x11_y51),
    .I1(x11_y58),
    .I2(x11_y51),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010100100101)
) lut_15_56 (
    .O(x15_y56),
    .I0(x13_y57),
    .I1(x12_y56),
    .I2(x12_y54),
    .I3(x13_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001110110000)
) lut_16_56 (
    .O(x16_y56),
    .I0(1'b0),
    .I1(x14_y54),
    .I2(x13_y57),
    .I3(x14_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011110011000)
) lut_17_56 (
    .O(x17_y56),
    .I0(x14_y57),
    .I1(1'b0),
    .I2(x15_y57),
    .I3(x15_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100000101010)
) lut_18_56 (
    .O(x18_y56),
    .I0(x15_y57),
    .I1(1'b0),
    .I2(x16_y54),
    .I3(x15_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110010111000)
) lut_19_56 (
    .O(x19_y56),
    .I0(x16_y58),
    .I1(x16_y60),
    .I2(x17_y55),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101111000011)
) lut_20_56 (
    .O(x20_y56),
    .I0(x17_y52),
    .I1(x18_y61),
    .I2(1'b0),
    .I3(x18_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010111011101)
) lut_21_56 (
    .O(x21_y56),
    .I0(x18_y56),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011010010010)
) lut_22_56 (
    .O(x22_y56),
    .I0(1'b0),
    .I1(x20_y57),
    .I2(x20_y54),
    .I3(x20_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111010001101)
) lut_23_56 (
    .O(x23_y56),
    .I0(x21_y57),
    .I1(x21_y52),
    .I2(x20_y56),
    .I3(x20_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001110000010)
) lut_24_56 (
    .O(x24_y56),
    .I0(x21_y55),
    .I1(1'b0),
    .I2(x22_y59),
    .I3(x22_y51)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001110101111)
) lut_25_56 (
    .O(x25_y56),
    .I0(1'b0),
    .I1(x22_y55),
    .I2(1'b0),
    .I3(x23_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011111101101)
) lut_26_56 (
    .O(x26_y56),
    .I0(x23_y59),
    .I1(x23_y59),
    .I2(1'b0),
    .I3(x24_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100101010010)
) lut_27_56 (
    .O(x27_y56),
    .I0(1'b0),
    .I1(x24_y60),
    .I2(x25_y54),
    .I3(x24_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110111100001)
) lut_28_56 (
    .O(x28_y56),
    .I0(x26_y59),
    .I1(1'b0),
    .I2(x26_y61),
    .I3(x26_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100001110101)
) lut_29_56 (
    .O(x29_y56),
    .I0(1'b0),
    .I1(x26_y58),
    .I2(1'b0),
    .I3(x26_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000001011110)
) lut_30_56 (
    .O(x30_y56),
    .I0(x27_y54),
    .I1(x28_y51),
    .I2(x28_y56),
    .I3(x27_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100001011111)
) lut_31_56 (
    .O(x31_y56),
    .I0(x29_y53),
    .I1(x28_y61),
    .I2(x29_y53),
    .I3(x28_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010011110100)
) lut_32_56 (
    .O(x32_y56),
    .I0(x29_y61),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x30_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001101010000)
) lut_33_56 (
    .O(x33_y56),
    .I0(x31_y57),
    .I1(1'b0),
    .I2(x31_y54),
    .I3(x31_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101101101000)
) lut_34_56 (
    .O(x34_y56),
    .I0(x32_y57),
    .I1(x31_y51),
    .I2(x32_y59),
    .I3(x31_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110001001001)
) lut_35_56 (
    .O(x35_y56),
    .I0(1'b0),
    .I1(x32_y54),
    .I2(x32_y52),
    .I3(x32_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101011101011)
) lut_36_56 (
    .O(x36_y56),
    .I0(x33_y53),
    .I1(1'b0),
    .I2(x34_y56),
    .I3(x34_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000100010100)
) lut_37_56 (
    .O(x37_y56),
    .I0(x34_y56),
    .I1(x35_y53),
    .I2(1'b0),
    .I3(x35_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011011010011)
) lut_38_56 (
    .O(x38_y56),
    .I0(x35_y61),
    .I1(x35_y56),
    .I2(x36_y59),
    .I3(x35_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010110111101)
) lut_39_56 (
    .O(x39_y56),
    .I0(1'b0),
    .I1(x36_y58),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101110111001)
) lut_40_56 (
    .O(x40_y56),
    .I0(x38_y53),
    .I1(x38_y55),
    .I2(x37_y53),
    .I3(x37_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110101100001)
) lut_41_56 (
    .O(x41_y56),
    .I0(x39_y54),
    .I1(x38_y53),
    .I2(1'b0),
    .I3(x38_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100011110101)
) lut_42_56 (
    .O(x42_y56),
    .I0(x39_y57),
    .I1(x40_y52),
    .I2(x39_y51),
    .I3(x40_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110001110000)
) lut_43_56 (
    .O(x43_y56),
    .I0(1'b0),
    .I1(x40_y53),
    .I2(x41_y59),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010100010100)
) lut_44_56 (
    .O(x44_y56),
    .I0(1'b0),
    .I1(x42_y61),
    .I2(x42_y54),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100110101010)
) lut_45_56 (
    .O(x45_y56),
    .I0(1'b0),
    .I1(x43_y54),
    .I2(x42_y55),
    .I3(x43_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111111100001)
) lut_46_56 (
    .O(x46_y56),
    .I0(1'b0),
    .I1(x43_y52),
    .I2(x44_y55),
    .I3(x43_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111011010011)
) lut_47_56 (
    .O(x47_y56),
    .I0(x44_y53),
    .I1(1'b0),
    .I2(x45_y56),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100110100000)
) lut_48_56 (
    .O(x48_y56),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x45_y60),
    .I3(x46_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100011101001)
) lut_49_56 (
    .O(x49_y56),
    .I0(x46_y53),
    .I1(x46_y51),
    .I2(x47_y53),
    .I3(x46_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100110110011)
) lut_50_56 (
    .O(x50_y56),
    .I0(x48_y53),
    .I1(x47_y54),
    .I2(x47_y60),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011000000000)
) lut_51_56 (
    .O(x51_y56),
    .I0(1'b0),
    .I1(x48_y57),
    .I2(x49_y51),
    .I3(x49_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110111000001)
) lut_52_56 (
    .O(x52_y56),
    .I0(x49_y61),
    .I1(x49_y61),
    .I2(x50_y58),
    .I3(x49_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000011010000)
) lut_53_56 (
    .O(x53_y56),
    .I0(x51_y61),
    .I1(x50_y59),
    .I2(x51_y61),
    .I3(x50_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110011100101)
) lut_54_56 (
    .O(x54_y56),
    .I0(x52_y57),
    .I1(x52_y54),
    .I2(x51_y53),
    .I3(x51_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100001011001)
) lut_55_56 (
    .O(x55_y56),
    .I0(x53_y57),
    .I1(x53_y57),
    .I2(x52_y52),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000111110000)
) lut_56_56 (
    .O(x56_y56),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x53_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011000000001)
) lut_57_56 (
    .O(x57_y56),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x55_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101011111001)
) lut_58_56 (
    .O(x58_y56),
    .I0(x56_y54),
    .I1(1'b0),
    .I2(x56_y60),
    .I3(x56_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010100110011)
) lut_59_56 (
    .O(x59_y56),
    .I0(x57_y59),
    .I1(x56_y54),
    .I2(1'b0),
    .I3(x57_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001001111011)
) lut_60_56 (
    .O(x60_y56),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x58_y57),
    .I3(x57_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011100100001)
) lut_61_56 (
    .O(x61_y56),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x59_y53),
    .I3(x59_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001100000011)
) lut_62_56 (
    .O(x62_y56),
    .I0(x60_y57),
    .I1(1'b0),
    .I2(x60_y61),
    .I3(x60_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011100001100)
) lut_0_57 (
    .O(x0_y57),
    .I0(1'b0),
    .I1(in2),
    .I2(in4),
    .I3(in1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001100111100)
) lut_1_57 (
    .O(x1_y57),
    .I0(in9),
    .I1(in1),
    .I2(in9),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010100101100)
) lut_2_57 (
    .O(x2_y57),
    .I0(in7),
    .I1(in2),
    .I2(in5),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000110110110)
) lut_3_57 (
    .O(x3_y57),
    .I0(1'b0),
    .I1(x1_y52),
    .I2(in5),
    .I3(x1_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111101011010)
) lut_4_57 (
    .O(x4_y57),
    .I0(x2_y56),
    .I1(1'b0),
    .I2(x2_y55),
    .I3(x2_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111110100101)
) lut_5_57 (
    .O(x5_y57),
    .I0(1'b0),
    .I1(x2_y59),
    .I2(x2_y60),
    .I3(x3_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000110100001)
) lut_6_57 (
    .O(x6_y57),
    .I0(x4_y53),
    .I1(x4_y61),
    .I2(1'b0),
    .I3(x4_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110000101101)
) lut_7_57 (
    .O(x7_y57),
    .I0(x5_y62),
    .I1(x5_y59),
    .I2(x5_y54),
    .I3(x5_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001100010101)
) lut_8_57 (
    .O(x8_y57),
    .I0(x5_y55),
    .I1(x5_y53),
    .I2(x5_y53),
    .I3(x6_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000001101110)
) lut_9_57 (
    .O(x9_y57),
    .I0(x6_y59),
    .I1(1'b0),
    .I2(x5_y53),
    .I3(x6_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110100111000)
) lut_10_57 (
    .O(x10_y57),
    .I0(x8_y61),
    .I1(x7_y57),
    .I2(x8_y57),
    .I3(x7_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111000100111)
) lut_11_57 (
    .O(x11_y57),
    .I0(x8_y57),
    .I1(1'b0),
    .I2(x8_y57),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110100100001)
) lut_12_57 (
    .O(x12_y57),
    .I0(x10_y61),
    .I1(x9_y55),
    .I2(x10_y61),
    .I3(x10_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111111100010)
) lut_13_57 (
    .O(x13_y57),
    .I0(x10_y58),
    .I1(x11_y56),
    .I2(x10_y55),
    .I3(x11_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000111111100)
) lut_14_57 (
    .O(x14_y57),
    .I0(1'b0),
    .I1(x12_y59),
    .I2(x12_y58),
    .I3(x11_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000100000100)
) lut_15_57 (
    .O(x15_y57),
    .I0(x13_y52),
    .I1(x12_y61),
    .I2(x13_y52),
    .I3(x12_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000010011110)
) lut_16_57 (
    .O(x16_y57),
    .I0(x13_y61),
    .I1(1'b0),
    .I2(x14_y61),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010110110011)
) lut_17_57 (
    .O(x17_y57),
    .I0(1'b0),
    .I1(x15_y57),
    .I2(x15_y55),
    .I3(x14_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100001001100)
) lut_18_57 (
    .O(x18_y57),
    .I0(x15_y56),
    .I1(x15_y56),
    .I2(x15_y57),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110111000001)
) lut_19_57 (
    .O(x19_y57),
    .I0(x16_y55),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x16_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011111011111)
) lut_20_57 (
    .O(x20_y57),
    .I0(1'b0),
    .I1(x18_y54),
    .I2(x17_y59),
    .I3(x17_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000011000010)
) lut_21_57 (
    .O(x21_y57),
    .I0(x19_y61),
    .I1(1'b0),
    .I2(x19_y53),
    .I3(x18_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110100011000)
) lut_22_57 (
    .O(x22_y57),
    .I0(x20_y54),
    .I1(x20_y58),
    .I2(x20_y61),
    .I3(x20_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001000100110)
) lut_23_57 (
    .O(x23_y57),
    .I0(x21_y53),
    .I1(1'b0),
    .I2(x20_y61),
    .I3(x21_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011000101010)
) lut_24_57 (
    .O(x24_y57),
    .I0(x21_y56),
    .I1(x22_y56),
    .I2(1'b0),
    .I3(x21_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101001010101)
) lut_25_57 (
    .O(x25_y57),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x23_y60),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001001010001)
) lut_26_57 (
    .O(x26_y57),
    .I0(1'b0),
    .I1(x24_y61),
    .I2(x23_y61),
    .I3(x24_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111011001000)
) lut_27_57 (
    .O(x27_y57),
    .I0(x25_y56),
    .I1(x24_y55),
    .I2(x25_y57),
    .I3(x24_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001000111110)
) lut_28_57 (
    .O(x28_y57),
    .I0(x25_y58),
    .I1(x25_y53),
    .I2(x26_y55),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111101011100)
) lut_29_57 (
    .O(x29_y57),
    .I0(x26_y57),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x26_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001010001100)
) lut_30_57 (
    .O(x30_y57),
    .I0(x27_y61),
    .I1(x27_y59),
    .I2(x27_y60),
    .I3(x27_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101100000101)
) lut_31_57 (
    .O(x31_y57),
    .I0(1'b0),
    .I1(x29_y53),
    .I2(x28_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011010011110)
) lut_32_57 (
    .O(x32_y57),
    .I0(x29_y62),
    .I1(x29_y62),
    .I2(x30_y61),
    .I3(x29_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001100001100)
) lut_33_57 (
    .O(x33_y57),
    .I0(x30_y56),
    .I1(x31_y60),
    .I2(x30_y57),
    .I3(x30_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000011111001)
) lut_34_57 (
    .O(x34_y57),
    .I0(x32_y60),
    .I1(x31_y62),
    .I2(x31_y55),
    .I3(x32_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101000100000)
) lut_35_57 (
    .O(x35_y57),
    .I0(x32_y57),
    .I1(x33_y55),
    .I2(x33_y52),
    .I3(x33_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000000100010)
) lut_36_57 (
    .O(x36_y57),
    .I0(x33_y59),
    .I1(x33_y53),
    .I2(x33_y57),
    .I3(x33_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101010001101)
) lut_37_57 (
    .O(x37_y57),
    .I0(1'b0),
    .I1(x34_y56),
    .I2(x34_y52),
    .I3(x34_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100000010000)
) lut_38_57 (
    .O(x38_y57),
    .I0(x35_y62),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100010111111)
) lut_39_57 (
    .O(x39_y57),
    .I0(x37_y61),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x36_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010100010101)
) lut_40_57 (
    .O(x40_y57),
    .I0(x37_y55),
    .I1(x38_y58),
    .I2(x37_y59),
    .I3(x37_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110100011000)
) lut_41_57 (
    .O(x41_y57),
    .I0(x39_y54),
    .I1(x38_y61),
    .I2(x39_y62),
    .I3(x39_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111111110101)
) lut_42_57 (
    .O(x42_y57),
    .I0(x39_y54),
    .I1(x39_y61),
    .I2(x40_y52),
    .I3(x39_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001101111010)
) lut_43_57 (
    .O(x43_y57),
    .I0(x40_y56),
    .I1(x40_y60),
    .I2(1'b0),
    .I3(x40_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101000111101)
) lut_44_57 (
    .O(x44_y57),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x41_y59),
    .I3(x41_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000100010001)
) lut_45_57 (
    .O(x45_y57),
    .I0(x42_y60),
    .I1(x43_y54),
    .I2(x42_y53),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010010001110)
) lut_46_57 (
    .O(x46_y57),
    .I0(x43_y56),
    .I1(x44_y55),
    .I2(1'b0),
    .I3(x43_y53)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100000011010)
) lut_47_57 (
    .O(x47_y57),
    .I0(x45_y61),
    .I1(x44_y56),
    .I2(x44_y58),
    .I3(x45_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001100011110)
) lut_48_57 (
    .O(x48_y57),
    .I0(x46_y60),
    .I1(x46_y61),
    .I2(x46_y56),
    .I3(x45_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011110111110)
) lut_49_57 (
    .O(x49_y57),
    .I0(x47_y62),
    .I1(x47_y62),
    .I2(1'b0),
    .I3(x47_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000100111000)
) lut_50_57 (
    .O(x50_y57),
    .I0(x48_y52),
    .I1(x48_y58),
    .I2(x47_y57),
    .I3(x48_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111110010001)
) lut_51_57 (
    .O(x51_y57),
    .I0(x49_y56),
    .I1(x49_y58),
    .I2(1'b0),
    .I3(x49_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101100101001)
) lut_52_57 (
    .O(x52_y57),
    .I0(x50_y55),
    .I1(x49_y59),
    .I2(x49_y59),
    .I3(x49_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011010101001)
) lut_53_57 (
    .O(x53_y57),
    .I0(1'b0),
    .I1(x51_y54),
    .I2(x51_y61),
    .I3(x50_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010100101010)
) lut_54_57 (
    .O(x54_y57),
    .I0(x51_y58),
    .I1(x51_y59),
    .I2(x52_y56),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110111001110)
) lut_55_57 (
    .O(x55_y57),
    .I0(x53_y52),
    .I1(x52_y56),
    .I2(x52_y52),
    .I3(x53_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100001001011)
) lut_56_57 (
    .O(x56_y57),
    .I0(x54_y58),
    .I1(x53_y56),
    .I2(x53_y59),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001110001110)
) lut_57_57 (
    .O(x57_y57),
    .I0(x55_y62),
    .I1(x55_y58),
    .I2(x55_y55),
    .I3(x54_y52)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111101011011)
) lut_58_57 (
    .O(x58_y57),
    .I0(1'b0),
    .I1(x55_y56),
    .I2(x55_y55),
    .I3(x55_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100100011100)
) lut_59_57 (
    .O(x59_y57),
    .I0(1'b0),
    .I1(x57_y54),
    .I2(1'b0),
    .I3(x56_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101101110101)
) lut_60_57 (
    .O(x60_y57),
    .I0(x58_y58),
    .I1(x57_y55),
    .I2(x58_y58),
    .I3(x57_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101100100110)
) lut_61_57 (
    .O(x61_y57),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101101101100)
) lut_62_57 (
    .O(x62_y57),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x59_y59),
    .I3(x59_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100101101100)
) lut_0_58 (
    .O(x0_y58),
    .I0(1'b0),
    .I1(in8),
    .I2(in7),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111111000101)
) lut_1_58 (
    .O(x1_y58),
    .I0(in4),
    .I1(in9),
    .I2(in7),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100010010000)
) lut_2_58 (
    .O(x2_y58),
    .I0(in6),
    .I1(in3),
    .I2(in2),
    .I3(in4)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101100100011)
) lut_3_58 (
    .O(x3_y58),
    .I0(x1_y55),
    .I1(x1_y55),
    .I2(x1_y57),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101110101000)
) lut_4_58 (
    .O(x4_y58),
    .I0(x2_y59),
    .I1(x1_y56),
    .I2(x2_y59),
    .I3(x2_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011000001010)
) lut_5_58 (
    .O(x5_y58),
    .I0(x2_y55),
    .I1(1'b0),
    .I2(x3_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011100100111)
) lut_6_58 (
    .O(x6_y58),
    .I0(x3_y58),
    .I1(x4_y58),
    .I2(x4_y54),
    .I3(x4_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100011011100)
) lut_7_58 (
    .O(x7_y58),
    .I0(x5_y53),
    .I1(x4_y54),
    .I2(x4_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001110001110)
) lut_8_58 (
    .O(x8_y58),
    .I0(x5_y56),
    .I1(x5_y60),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101110100000)
) lut_9_58 (
    .O(x9_y58),
    .I0(x6_y57),
    .I1(x7_y62),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011010001100)
) lut_10_58 (
    .O(x10_y58),
    .I0(x8_y60),
    .I1(1'b0),
    .I2(x7_y57),
    .I3(x7_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100111111111)
) lut_11_58 (
    .O(x11_y58),
    .I0(1'b0),
    .I1(x9_y53),
    .I2(x9_y62),
    .I3(x8_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101000111010)
) lut_12_58 (
    .O(x12_y58),
    .I0(x10_y53),
    .I1(x10_y56),
    .I2(x10_y55),
    .I3(x10_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110000010010)
) lut_13_58 (
    .O(x13_y58),
    .I0(x10_y57),
    .I1(1'b0),
    .I2(x10_y53),
    .I3(x10_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111110001111)
) lut_14_58 (
    .O(x14_y58),
    .I0(1'b0),
    .I1(x12_y55),
    .I2(1'b0),
    .I3(x12_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111011011111)
) lut_15_58 (
    .O(x15_y58),
    .I0(x13_y56),
    .I1(x13_y55),
    .I2(x12_y59),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110110101111)
) lut_16_58 (
    .O(x16_y58),
    .I0(1'b0),
    .I1(x13_y59),
    .I2(x13_y57),
    .I3(x13_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000000000011)
) lut_17_58 (
    .O(x17_y58),
    .I0(x15_y58),
    .I1(x15_y53),
    .I2(x14_y60),
    .I3(x15_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001101010101)
) lut_18_58 (
    .O(x18_y58),
    .I0(x16_y53),
    .I1(x16_y61),
    .I2(x15_y55),
    .I3(x16_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011010010011)
) lut_19_58 (
    .O(x19_y58),
    .I0(x16_y60),
    .I1(x17_y62),
    .I2(x17_y59),
    .I3(x17_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110000100011)
) lut_20_58 (
    .O(x20_y58),
    .I0(x18_y60),
    .I1(1'b0),
    .I2(x17_y62),
    .I3(x18_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111101111011)
) lut_21_58 (
    .O(x21_y58),
    .I0(x18_y61),
    .I1(x18_y55),
    .I2(x19_y55),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011000101111)
) lut_22_58 (
    .O(x22_y58),
    .I0(x19_y58),
    .I1(x19_y61),
    .I2(x19_y61),
    .I3(x19_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011100001100)
) lut_23_58 (
    .O(x23_y58),
    .I0(1'b0),
    .I1(x21_y53),
    .I2(x20_y61),
    .I3(x20_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010011111111)
) lut_24_58 (
    .O(x24_y58),
    .I0(x21_y54),
    .I1(1'b0),
    .I2(x22_y61),
    .I3(x21_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011100001001)
) lut_25_58 (
    .O(x25_y58),
    .I0(x23_y54),
    .I1(x22_y54),
    .I2(x23_y55),
    .I3(x22_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011111111101)
) lut_26_58 (
    .O(x26_y58),
    .I0(x24_y60),
    .I1(x23_y62),
    .I2(1'b0),
    .I3(x24_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111111101010)
) lut_27_58 (
    .O(x27_y58),
    .I0(x25_y62),
    .I1(x25_y54),
    .I2(x25_y53),
    .I3(x25_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000011101001)
) lut_28_58 (
    .O(x28_y58),
    .I0(x26_y55),
    .I1(x25_y61),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110010011101)
) lut_29_58 (
    .O(x29_y58),
    .I0(1'b0),
    .I1(x26_y58),
    .I2(x27_y61),
    .I3(x27_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101111010010)
) lut_30_58 (
    .O(x30_y58),
    .I0(x27_y54),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111011011100)
) lut_31_58 (
    .O(x31_y58),
    .I0(x29_y53),
    .I1(1'b0),
    .I2(x29_y53),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011101001110)
) lut_32_58 (
    .O(x32_y58),
    .I0(1'b0),
    .I1(x29_y60),
    .I2(x29_y54),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000000000000)
) lut_33_58 (
    .O(x33_y58),
    .I0(x30_y54),
    .I1(x30_y59),
    .I2(1'b0),
    .I3(x30_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110110111011)
) lut_34_58 (
    .O(x34_y58),
    .I0(x31_y53),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101111000000)
) lut_35_58 (
    .O(x35_y58),
    .I0(1'b0),
    .I1(x33_y57),
    .I2(1'b0),
    .I3(x33_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010010000111)
) lut_36_58 (
    .O(x36_y58),
    .I0(x33_y59),
    .I1(x33_y55),
    .I2(x33_y53),
    .I3(x34_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000011111010)
) lut_37_58 (
    .O(x37_y58),
    .I0(1'b0),
    .I1(x34_y56),
    .I2(x35_y60),
    .I3(x35_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001111100101)
) lut_38_58 (
    .O(x38_y58),
    .I0(x36_y58),
    .I1(1'b0),
    .I2(x36_y53),
    .I3(x35_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111001110111)
) lut_39_58 (
    .O(x39_y58),
    .I0(x37_y62),
    .I1(1'b0),
    .I2(x36_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110100110110)
) lut_40_58 (
    .O(x40_y58),
    .I0(x37_y62),
    .I1(x38_y55),
    .I2(1'b0),
    .I3(x38_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111000110011)
) lut_41_58 (
    .O(x41_y58),
    .I0(x39_y59),
    .I1(x38_y59),
    .I2(1'b0),
    .I3(x39_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011001000010)
) lut_42_58 (
    .O(x42_y58),
    .I0(x39_y62),
    .I1(1'b0),
    .I2(x39_y58),
    .I3(x39_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110110010011)
) lut_43_58 (
    .O(x43_y58),
    .I0(x40_y53),
    .I1(x41_y53),
    .I2(x41_y62),
    .I3(x41_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010001011111)
) lut_44_58 (
    .O(x44_y58),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100011001011)
) lut_45_58 (
    .O(x45_y58),
    .I0(x42_y61),
    .I1(x43_y57),
    .I2(x42_y61),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001011001010)
) lut_46_58 (
    .O(x46_y58),
    .I0(x44_y55),
    .I1(x43_y59),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100100000100)
) lut_47_58 (
    .O(x47_y58),
    .I0(x44_y62),
    .I1(1'b0),
    .I2(x45_y62),
    .I3(x45_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101000101111)
) lut_48_58 (
    .O(x48_y58),
    .I0(x45_y54),
    .I1(x46_y58),
    .I2(1'b0),
    .I3(x46_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110000100011)
) lut_49_58 (
    .O(x49_y58),
    .I0(x46_y61),
    .I1(1'b0),
    .I2(x46_y61),
    .I3(x46_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101110010011)
) lut_50_58 (
    .O(x50_y58),
    .I0(x48_y56),
    .I1(x48_y61),
    .I2(x47_y58),
    .I3(x48_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110010101000)
) lut_51_58 (
    .O(x51_y58),
    .I0(x48_y62),
    .I1(1'b0),
    .I2(x49_y55),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010011111101)
) lut_52_58 (
    .O(x52_y58),
    .I0(x50_y55),
    .I1(x49_y58),
    .I2(x50_y56),
    .I3(x50_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001100101000)
) lut_53_58 (
    .O(x53_y58),
    .I0(x51_y61),
    .I1(1'b0),
    .I2(x50_y57),
    .I3(x50_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101101001001)
) lut_54_58 (
    .O(x54_y58),
    .I0(x52_y55),
    .I1(x52_y58),
    .I2(x51_y57),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001111001111)
) lut_55_58 (
    .O(x55_y58),
    .I0(x53_y58),
    .I1(x53_y55),
    .I2(x53_y58),
    .I3(x53_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000111001100)
) lut_56_58 (
    .O(x56_y58),
    .I0(x54_y55),
    .I1(x53_y56),
    .I2(x53_y53),
    .I3(x54_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101010001111)
) lut_57_58 (
    .O(x57_y58),
    .I0(x55_y53),
    .I1(1'b0),
    .I2(x54_y55),
    .I3(x54_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011110000010)
) lut_58_58 (
    .O(x58_y58),
    .I0(x56_y55),
    .I1(x55_y55),
    .I2(1'b0),
    .I3(x55_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100101011000)
) lut_59_58 (
    .O(x59_y58),
    .I0(x56_y62),
    .I1(1'b0),
    .I2(x56_y62),
    .I3(x56_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001100101111)
) lut_60_58 (
    .O(x60_y58),
    .I0(x58_y62),
    .I1(x58_y58),
    .I2(x57_y57),
    .I3(x58_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111111000001)
) lut_61_58 (
    .O(x61_y58),
    .I0(x59_y62),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x58_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101011010100)
) lut_62_58 (
    .O(x62_y58),
    .I0(x60_y53),
    .I1(1'b0),
    .I2(x60_y60),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100011011100)
) lut_0_59 (
    .O(x0_y59),
    .I0(1'b0),
    .I1(in8),
    .I2(in1),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001101111101)
) lut_1_59 (
    .O(x1_y59),
    .I0(in2),
    .I1(1'b0),
    .I2(in6),
    .I3(in7)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011011010110)
) lut_2_59 (
    .O(x2_y59),
    .I0(in7),
    .I1(1'b0),
    .I2(in7),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111000111111)
) lut_3_59 (
    .O(x3_y59),
    .I0(in2),
    .I1(x1_y54),
    .I2(1'b0),
    .I3(x1_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010110110000)
) lut_4_59 (
    .O(x4_y59),
    .I0(x2_y61),
    .I1(x1_y60),
    .I2(1'b0),
    .I3(x1_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000010010110)
) lut_5_59 (
    .O(x5_y59),
    .I0(x2_y61),
    .I1(x3_y60),
    .I2(x3_y61),
    .I3(x2_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010010101101)
) lut_6_59 (
    .O(x6_y59),
    .I0(x3_y62),
    .I1(x3_y58),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101001001101)
) lut_7_59 (
    .O(x7_y59),
    .I0(x5_y56),
    .I1(x4_y58),
    .I2(1'b0),
    .I3(x4_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010010111110)
) lut_8_59 (
    .O(x8_y59),
    .I0(x6_y54),
    .I1(x5_y54),
    .I2(x6_y55),
    .I3(x5_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011011111010)
) lut_9_59 (
    .O(x9_y59),
    .I0(x6_y62),
    .I1(1'b0),
    .I2(x6_y55),
    .I3(x5_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100001000010)
) lut_10_59 (
    .O(x10_y59),
    .I0(x7_y56),
    .I1(x8_y62),
    .I2(x7_y58),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111101011100)
) lut_11_59 (
    .O(x11_y59),
    .I0(x8_y62),
    .I1(x8_y57),
    .I2(x9_y58),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111001101101)
) lut_12_59 (
    .O(x12_y59),
    .I0(x9_y62),
    .I1(x9_y62),
    .I2(x9_y58),
    .I3(x10_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010110101101)
) lut_13_59 (
    .O(x13_y59),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x11_y59),
    .I3(x10_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010010010000)
) lut_14_59 (
    .O(x14_y59),
    .I0(x11_y58),
    .I1(1'b0),
    .I2(x11_y57),
    .I3(x12_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100000001010)
) lut_15_59 (
    .O(x15_y59),
    .I0(x13_y57),
    .I1(x12_y57),
    .I2(x13_y54),
    .I3(x12_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001001000101)
) lut_16_59 (
    .O(x16_y59),
    .I0(x14_y55),
    .I1(x14_y59),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110011001110)
) lut_17_59 (
    .O(x17_y59),
    .I0(x15_y59),
    .I1(1'b0),
    .I2(x14_y57),
    .I3(x15_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000100110111)
) lut_18_59 (
    .O(x18_y59),
    .I0(x16_y59),
    .I1(x16_y62),
    .I2(x16_y58),
    .I3(x15_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101011000000)
) lut_19_59 (
    .O(x19_y59),
    .I0(1'b0),
    .I1(x16_y54),
    .I2(x17_y57),
    .I3(x16_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100000110001)
) lut_20_59 (
    .O(x20_y59),
    .I0(x18_y62),
    .I1(x17_y56),
    .I2(x18_y62),
    .I3(x18_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110100010100)
) lut_21_59 (
    .O(x21_y59),
    .I0(1'b0),
    .I1(x19_y60),
    .I2(x18_y56),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001010000111)
) lut_22_59 (
    .O(x22_y59),
    .I0(x19_y54),
    .I1(x20_y62),
    .I2(x19_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011000100010)
) lut_23_59 (
    .O(x23_y59),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x21_y62),
    .I3(x20_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100110111100)
) lut_24_59 (
    .O(x24_y59),
    .I0(x22_y60),
    .I1(x21_y55),
    .I2(1'b0),
    .I3(x22_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101111100100)
) lut_25_59 (
    .O(x25_y59),
    .I0(x22_y62),
    .I1(x22_y59),
    .I2(x22_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000000111111)
) lut_26_59 (
    .O(x26_y59),
    .I0(x23_y58),
    .I1(1'b0),
    .I2(x24_y55),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100101010011)
) lut_27_59 (
    .O(x27_y59),
    .I0(x24_y54),
    .I1(x25_y60),
    .I2(1'b0),
    .I3(x24_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110101100101)
) lut_28_59 (
    .O(x28_y59),
    .I0(1'b0),
    .I1(x25_y62),
    .I2(x26_y55),
    .I3(x25_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000000010000)
) lut_29_59 (
    .O(x29_y59),
    .I0(x27_y60),
    .I1(x27_y60),
    .I2(x26_y58),
    .I3(x26_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110111110001)
) lut_30_59 (
    .O(x30_y59),
    .I0(x28_y62),
    .I1(x28_y56),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001101011100)
) lut_31_59 (
    .O(x31_y59),
    .I0(x29_y55),
    .I1(x28_y62),
    .I2(x29_y62),
    .I3(x28_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100000101001)
) lut_32_59 (
    .O(x32_y59),
    .I0(x29_y56),
    .I1(x30_y57),
    .I2(x30_y59),
    .I3(x29_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100000100001)
) lut_33_59 (
    .O(x33_y59),
    .I0(x30_y61),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001001110001)
) lut_34_59 (
    .O(x34_y59),
    .I0(1'b0),
    .I1(x31_y61),
    .I2(x31_y57),
    .I3(x31_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110100101101)
) lut_35_59 (
    .O(x35_y59),
    .I0(x33_y62),
    .I1(x33_y55),
    .I2(x32_y57),
    .I3(x32_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000000000001)
) lut_36_59 (
    .O(x36_y59),
    .I0(x33_y62),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x34_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010100010011)
) lut_37_59 (
    .O(x37_y59),
    .I0(x35_y58),
    .I1(x34_y55),
    .I2(x34_y54),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110100000001)
) lut_38_59 (
    .O(x38_y59),
    .I0(x36_y55),
    .I1(1'b0),
    .I2(x36_y58),
    .I3(x35_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011111110110)
) lut_39_59 (
    .O(x39_y59),
    .I0(1'b0),
    .I1(x37_y56),
    .I2(x37_y54),
    .I3(x37_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110101110111)
) lut_40_59 (
    .O(x40_y59),
    .I0(x38_y62),
    .I1(x37_y54),
    .I2(1'b0),
    .I3(x38_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010101001011)
) lut_41_59 (
    .O(x41_y59),
    .I0(x38_y62),
    .I1(x38_y60),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101011110111)
) lut_42_59 (
    .O(x42_y59),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x40_y57),
    .I3(x40_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011000110100)
) lut_43_59 (
    .O(x43_y59),
    .I0(x41_y62),
    .I1(x40_y61),
    .I2(x40_y62),
    .I3(x41_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011001001101)
) lut_44_59 (
    .O(x44_y59),
    .I0(x41_y62),
    .I1(x42_y60),
    .I2(x42_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101001010000)
) lut_45_59 (
    .O(x45_y59),
    .I0(1'b0),
    .I1(x42_y56),
    .I2(1'b0),
    .I3(x43_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100001101001)
) lut_46_59 (
    .O(x46_y59),
    .I0(1'b0),
    .I1(x44_y62),
    .I2(x44_y57),
    .I3(x44_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110010001110)
) lut_47_59 (
    .O(x47_y59),
    .I0(1'b0),
    .I1(x45_y56),
    .I2(x44_y59),
    .I3(x45_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100111000110)
) lut_48_59 (
    .O(x48_y59),
    .I0(x46_y57),
    .I1(x46_y61),
    .I2(x45_y60),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110111001111)
) lut_49_59 (
    .O(x49_y59),
    .I0(x46_y57),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100110110011)
) lut_50_59 (
    .O(x50_y59),
    .I0(x47_y62),
    .I1(x47_y57),
    .I2(x48_y54),
    .I3(x48_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010011001001)
) lut_51_59 (
    .O(x51_y59),
    .I0(x48_y62),
    .I1(x49_y57),
    .I2(x48_y56),
    .I3(x49_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011011110111)
) lut_52_59 (
    .O(x52_y59),
    .I0(x50_y55),
    .I1(x49_y56),
    .I2(x50_y60),
    .I3(x49_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011111011010)
) lut_53_59 (
    .O(x53_y59),
    .I0(x50_y62),
    .I1(1'b0),
    .I2(x51_y55),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101001100001)
) lut_54_59 (
    .O(x54_y59),
    .I0(1'b0),
    .I1(x52_y62),
    .I2(x51_y60),
    .I3(x52_y54)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010110111011)
) lut_55_59 (
    .O(x55_y59),
    .I0(1'b0),
    .I1(x53_y62),
    .I2(1'b0),
    .I3(x53_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010100000100)
) lut_56_59 (
    .O(x56_y59),
    .I0(x53_y57),
    .I1(x54_y62),
    .I2(1'b0),
    .I3(x53_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111110110110)
) lut_57_59 (
    .O(x57_y59),
    .I0(x55_y62),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001010111110)
) lut_58_59 (
    .O(x58_y59),
    .I0(x55_y58),
    .I1(x55_y62),
    .I2(x56_y60),
    .I3(x55_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101110110101)
) lut_59_59 (
    .O(x59_y59),
    .I0(x57_y62),
    .I1(x57_y54),
    .I2(x57_y54),
    .I3(x57_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001001110100)
) lut_60_59 (
    .O(x60_y59),
    .I0(x57_y55),
    .I1(1'b0),
    .I2(x58_y54),
    .I3(x57_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100001111010)
) lut_61_59 (
    .O(x61_y59),
    .I0(x59_y61),
    .I1(x59_y62),
    .I2(x59_y55),
    .I3(x58_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011110100110)
) lut_62_59 (
    .O(x62_y59),
    .I0(1'b0),
    .I1(x60_y59),
    .I2(x59_y55),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110001111111)
) lut_0_60 (
    .O(x0_y60),
    .I0(in1),
    .I1(in2),
    .I2(1'b0),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111100111000)
) lut_1_60 (
    .O(x1_y60),
    .I0(in2),
    .I1(in2),
    .I2(in6),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010101010110)
) lut_2_60 (
    .O(x2_y60),
    .I0(in2),
    .I1(in9),
    .I2(in2),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101000010111)
) lut_3_60 (
    .O(x3_y60),
    .I0(in8),
    .I1(1'b0),
    .I2(x1_y55),
    .I3(x1_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100011111110)
) lut_4_60 (
    .O(x4_y60),
    .I0(1'b0),
    .I1(x2_y62),
    .I2(x2_y57),
    .I3(x2_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001000101111)
) lut_5_60 (
    .O(x5_y60),
    .I0(x2_y62),
    .I1(x2_y61),
    .I2(1'b0),
    .I3(x2_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000011101011)
) lut_6_60 (
    .O(x6_y60),
    .I0(x3_y62),
    .I1(x3_y56),
    .I2(x4_y56),
    .I3(x4_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110101000011)
) lut_7_60 (
    .O(x7_y60),
    .I0(x5_y61),
    .I1(x5_y60),
    .I2(x4_y57),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000100101010)
) lut_8_60 (
    .O(x8_y60),
    .I0(x6_y62),
    .I1(1'b0),
    .I2(x5_y58),
    .I3(x6_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100001000011)
) lut_9_60 (
    .O(x9_y60),
    .I0(x7_y56),
    .I1(1'b0),
    .I2(x5_y58),
    .I3(x6_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111001010100)
) lut_10_60 (
    .O(x10_y60),
    .I0(x8_y62),
    .I1(x7_y62),
    .I2(x8_y56),
    .I3(x7_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111110111001)
) lut_11_60 (
    .O(x11_y60),
    .I0(1'b0),
    .I1(x9_y61),
    .I2(x9_y57),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010110101111)
) lut_12_60 (
    .O(x12_y60),
    .I0(1'b0),
    .I1(x9_y62),
    .I2(x10_y61),
    .I3(x9_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110010001111)
) lut_13_60 (
    .O(x13_y60),
    .I0(x10_y56),
    .I1(x11_y62),
    .I2(x11_y58),
    .I3(x10_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001011110101)
) lut_14_60 (
    .O(x14_y60),
    .I0(x11_y60),
    .I1(x11_y62),
    .I2(1'b0),
    .I3(x11_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111111101100)
) lut_15_60 (
    .O(x15_y60),
    .I0(x13_y60),
    .I1(x12_y62),
    .I2(x12_y57),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001101010101)
) lut_16_60 (
    .O(x16_y60),
    .I0(x14_y59),
    .I1(1'b0),
    .I2(x14_y55),
    .I3(x14_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110100010001)
) lut_17_60 (
    .O(x17_y60),
    .I0(x14_y58),
    .I1(x14_y62),
    .I2(1'b0),
    .I3(x15_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011101110110)
) lut_18_60 (
    .O(x18_y60),
    .I0(x16_y62),
    .I1(x16_y57),
    .I2(x15_y55),
    .I3(x16_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101100101011)
) lut_19_60 (
    .O(x19_y60),
    .I0(x16_y58),
    .I1(x16_y62),
    .I2(x17_y60),
    .I3(x16_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111100010011)
) lut_20_60 (
    .O(x20_y60),
    .I0(x18_y56),
    .I1(x17_y62),
    .I2(x18_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010001011110)
) lut_21_60 (
    .O(x21_y60),
    .I0(1'b0),
    .I1(x18_y59),
    .I2(x18_y59),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001101011001)
) lut_22_60 (
    .O(x22_y60),
    .I0(x19_y60),
    .I1(x19_y55),
    .I2(x20_y62),
    .I3(x20_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110011010010)
) lut_23_60 (
    .O(x23_y60),
    .I0(x21_y55),
    .I1(x20_y60),
    .I2(1'b0),
    .I3(x20_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010100001001)
) lut_24_60 (
    .O(x24_y60),
    .I0(x22_y61),
    .I1(1'b0),
    .I2(x21_y57),
    .I3(x21_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110101011001)
) lut_25_60 (
    .O(x25_y60),
    .I0(1'b0),
    .I1(x22_y59),
    .I2(1'b0),
    .I3(x22_y55)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011110010001)
) lut_26_60 (
    .O(x26_y60),
    .I0(1'b0),
    .I1(x24_y59),
    .I2(x23_y56),
    .I3(x23_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100001100111)
) lut_27_60 (
    .O(x27_y60),
    .I0(1'b0),
    .I1(x24_y62),
    .I2(x24_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100001100011)
) lut_28_60 (
    .O(x28_y60),
    .I0(1'b0),
    .I1(x26_y60),
    .I2(x26_y59),
    .I3(x25_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000010001110)
) lut_29_60 (
    .O(x29_y60),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x26_y62),
    .I3(x26_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010010000100)
) lut_30_60 (
    .O(x30_y60),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x28_y60),
    .I3(x28_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010001011101)
) lut_31_60 (
    .O(x31_y60),
    .I0(x28_y62),
    .I1(x29_y58),
    .I2(x28_y62),
    .I3(x28_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011101001100)
) lut_32_60 (
    .O(x32_y60),
    .I0(x30_y59),
    .I1(x29_y55),
    .I2(1'b0),
    .I3(x29_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000110101101)
) lut_33_60 (
    .O(x33_y60),
    .I0(x30_y60),
    .I1(x30_y56),
    .I2(x31_y58),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001010111011)
) lut_34_60 (
    .O(x34_y60),
    .I0(x31_y62),
    .I1(1'b0),
    .I2(x32_y58),
    .I3(x32_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110010100101)
) lut_35_60 (
    .O(x35_y60),
    .I0(x33_y62),
    .I1(x33_y62),
    .I2(x32_y62),
    .I3(x32_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110101000100)
) lut_36_60 (
    .O(x36_y60),
    .I0(x33_y62),
    .I1(x34_y62),
    .I2(x33_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000101000100)
) lut_37_60 (
    .O(x37_y60),
    .I0(1'b0),
    .I1(x35_y62),
    .I2(x34_y57),
    .I3(x34_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001100000010)
) lut_38_60 (
    .O(x38_y60),
    .I0(x35_y56),
    .I1(x36_y61),
    .I2(x35_y60),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011111010011)
) lut_39_60 (
    .O(x39_y60),
    .I0(1'b0),
    .I1(x37_y62),
    .I2(x36_y61),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100010110111)
) lut_40_60 (
    .O(x40_y60),
    .I0(x38_y62),
    .I1(x37_y57),
    .I2(x38_y61),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100010111100)
) lut_41_60 (
    .O(x41_y60),
    .I0(1'b0),
    .I1(x39_y59),
    .I2(x39_y55),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000111011111)
) lut_42_60 (
    .O(x42_y60),
    .I0(1'b0),
    .I1(x40_y60),
    .I2(x40_y60),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000011011010)
) lut_43_60 (
    .O(x43_y60),
    .I0(x40_y62),
    .I1(x41_y62),
    .I2(x41_y57),
    .I3(x40_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111100111101)
) lut_44_60 (
    .O(x44_y60),
    .I0(x42_y58),
    .I1(1'b0),
    .I2(x42_y62),
    .I3(x42_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100110100100)
) lut_45_60 (
    .O(x45_y60),
    .I0(x42_y60),
    .I1(1'b0),
    .I2(x43_y60),
    .I3(x42_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100101101010)
) lut_46_60 (
    .O(x46_y60),
    .I0(x43_y61),
    .I1(x43_y62),
    .I2(x44_y59),
    .I3(x43_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001101100101)
) lut_47_60 (
    .O(x47_y60),
    .I0(1'b0),
    .I1(x44_y59),
    .I2(x44_y59),
    .I3(x45_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100001010000)
) lut_48_60 (
    .O(x48_y60),
    .I0(x46_y62),
    .I1(x46_y62),
    .I2(1'b0),
    .I3(x46_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100011011100)
) lut_49_60 (
    .O(x49_y60),
    .I0(x46_y60),
    .I1(x46_y62),
    .I2(x47_y62),
    .I3(x46_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110001110010)
) lut_50_60 (
    .O(x50_y60),
    .I0(x47_y62),
    .I1(x47_y59),
    .I2(x47_y62),
    .I3(x48_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110011100111)
) lut_51_60 (
    .O(x51_y60),
    .I0(x49_y56),
    .I1(x49_y62),
    .I2(x48_y56),
    .I3(x48_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110010100011)
) lut_52_60 (
    .O(x52_y60),
    .I0(x49_y55),
    .I1(x50_y62),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011110100111)
) lut_53_60 (
    .O(x53_y60),
    .I0(x50_y55),
    .I1(x50_y59),
    .I2(x50_y62),
    .I3(x51_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101001000011)
) lut_54_60 (
    .O(x54_y60),
    .I0(x52_y62),
    .I1(1'b0),
    .I2(x52_y62),
    .I3(x52_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011011010101)
) lut_55_60 (
    .O(x55_y60),
    .I0(x52_y62),
    .I1(x53_y59),
    .I2(x52_y60),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100000011000)
) lut_56_60 (
    .O(x56_y60),
    .I0(x53_y56),
    .I1(x53_y55),
    .I2(1'b0),
    .I3(x53_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100011100011)
) lut_57_60 (
    .O(x57_y60),
    .I0(1'b0),
    .I1(x54_y62),
    .I2(x54_y58),
    .I3(x55_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100100011010)
) lut_58_60 (
    .O(x58_y60),
    .I0(1'b0),
    .I1(x56_y55),
    .I2(x55_y58),
    .I3(x55_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110011101101)
) lut_59_60 (
    .O(x59_y60),
    .I0(x56_y58),
    .I1(x57_y62),
    .I2(1'b0),
    .I3(x56_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011000000000)
) lut_60_60 (
    .O(x60_y60),
    .I0(1'b0),
    .I1(x57_y62),
    .I2(x57_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111011111011)
) lut_61_60 (
    .O(x61_y60),
    .I0(1'b0),
    .I1(x58_y62),
    .I2(x59_y56),
    .I3(x58_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001010100011)
) lut_62_60 (
    .O(x62_y60),
    .I0(x60_y57),
    .I1(x59_y62),
    .I2(x59_y57),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001101110111)
) lut_0_61 (
    .O(x0_y61),
    .I0(1'b0),
    .I1(in2),
    .I2(1'b0),
    .I3(in8)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100100111110)
) lut_1_61 (
    .O(x1_y61),
    .I0(in0),
    .I1(1'b0),
    .I2(in0),
    .I3(in1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100110110011)
) lut_2_61 (
    .O(x2_y61),
    .I0(in1),
    .I1(in1),
    .I2(in2),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111001010011)
) lut_3_61 (
    .O(x3_y61),
    .I0(1'b0),
    .I1(in9),
    .I2(1'b0),
    .I3(x1_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011111010000)
) lut_4_61 (
    .O(x4_y61),
    .I0(x2_y58),
    .I1(x2_y60),
    .I2(x1_y60),
    .I3(x1_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000101100010)
) lut_5_61 (
    .O(x5_y61),
    .I0(x2_y62),
    .I1(x3_y61),
    .I2(x2_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101101110110)
) lut_6_61 (
    .O(x6_y61),
    .I0(1'b0),
    .I1(x3_y62),
    .I2(1'b0),
    .I3(x3_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110110101000)
) lut_7_61 (
    .O(x7_y61),
    .I0(1'b0),
    .I1(x5_y60),
    .I2(x5_y59),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010001010101)
) lut_8_61 (
    .O(x8_y61),
    .I0(x5_y61),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001000010011)
) lut_9_61 (
    .O(x9_y61),
    .I0(x6_y59),
    .I1(x7_y62),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110001101111)
) lut_10_61 (
    .O(x10_y61),
    .I0(x7_y61),
    .I1(x8_y56),
    .I2(x8_y62),
    .I3(x8_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111110100100)
) lut_11_61 (
    .O(x11_y61),
    .I0(x8_y60),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x9_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100110001101)
) lut_12_61 (
    .O(x12_y61),
    .I0(1'b0),
    .I1(x10_y62),
    .I2(x10_y58),
    .I3(x9_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011100011011)
) lut_13_61 (
    .O(x13_y61),
    .I0(1'b0),
    .I1(x10_y61),
    .I2(x11_y62),
    .I3(x10_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011111110110)
) lut_14_61 (
    .O(x14_y61),
    .I0(x12_y59),
    .I1(x12_y62),
    .I2(x11_y62),
    .I3(x12_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000111100100)
) lut_15_61 (
    .O(x15_y61),
    .I0(x12_y62),
    .I1(1'b0),
    .I2(x13_y62),
    .I3(x12_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010000011011)
) lut_16_61 (
    .O(x16_y61),
    .I0(1'b0),
    .I1(x13_y60),
    .I2(1'b0),
    .I3(x13_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001111100100)
) lut_17_61 (
    .O(x17_y61),
    .I0(x15_y62),
    .I1(1'b0),
    .I2(x14_y61),
    .I3(x14_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111100110100)
) lut_18_61 (
    .O(x18_y61),
    .I0(x16_y62),
    .I1(x15_y61),
    .I2(x15_y61),
    .I3(x16_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111011011001)
) lut_19_61 (
    .O(x19_y61),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x17_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010110111010)
) lut_20_61 (
    .O(x20_y61),
    .I0(x18_y62),
    .I1(x17_y62),
    .I2(x17_y57),
    .I3(x17_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011110000010)
) lut_21_61 (
    .O(x21_y61),
    .I0(x18_y62),
    .I1(x18_y59),
    .I2(x18_y61),
    .I3(x19_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000110011000)
) lut_22_61 (
    .O(x22_y61),
    .I0(x19_y62),
    .I1(x19_y59),
    .I2(x19_y60),
    .I3(x20_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011011010100)
) lut_23_61 (
    .O(x23_y61),
    .I0(x21_y62),
    .I1(x21_y62),
    .I2(1'b0),
    .I3(x20_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111011100011)
) lut_24_61 (
    .O(x24_y61),
    .I0(x21_y56),
    .I1(x22_y61),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010111100110)
) lut_25_61 (
    .O(x25_y61),
    .I0(x22_y58),
    .I1(1'b0),
    .I2(x23_y62),
    .I3(x22_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011000001011)
) lut_26_61 (
    .O(x26_y61),
    .I0(x24_y62),
    .I1(x23_y62),
    .I2(x24_y60),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000111100101)
) lut_27_61 (
    .O(x27_y61),
    .I0(1'b0),
    .I1(x24_y60),
    .I2(x24_y60),
    .I3(x24_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010010101111)
) lut_28_61 (
    .O(x28_y61),
    .I0(x26_y60),
    .I1(x25_y56),
    .I2(x26_y62),
    .I3(x26_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111101110000)
) lut_29_61 (
    .O(x29_y61),
    .I0(1'b0),
    .I1(x27_y62),
    .I2(x27_y62),
    .I3(x27_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110111100011)
) lut_30_61 (
    .O(x30_y61),
    .I0(x28_y56),
    .I1(x28_y60),
    .I2(1'b0),
    .I3(x27_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110111111011)
) lut_31_61 (
    .O(x31_y61),
    .I0(1'b0),
    .I1(x29_y62),
    .I2(x28_y56),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000010100011)
) lut_32_61 (
    .O(x32_y61),
    .I0(x29_y62),
    .I1(x29_y56),
    .I2(x29_y62),
    .I3(x30_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101100110001)
) lut_33_61 (
    .O(x33_y61),
    .I0(x31_y60),
    .I1(x31_y58),
    .I2(x31_y57),
    .I3(x30_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000111010111)
) lut_34_61 (
    .O(x34_y61),
    .I0(x31_y56),
    .I1(x31_y62),
    .I2(1'b0),
    .I3(x32_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011110011001)
) lut_35_61 (
    .O(x35_y61),
    .I0(x33_y60),
    .I1(1'b0),
    .I2(x33_y56),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000100101111)
) lut_36_61 (
    .O(x36_y61),
    .I0(x34_y59),
    .I1(x34_y62),
    .I2(x33_y58),
    .I3(x34_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001100101010)
) lut_37_61 (
    .O(x37_y61),
    .I0(x34_y60),
    .I1(x35_y62),
    .I2(1'b0),
    .I3(x34_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011001010101)
) lut_38_61 (
    .O(x38_y61),
    .I0(x35_y62),
    .I1(x35_y59),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011000001011)
) lut_39_61 (
    .O(x39_y61),
    .I0(x37_y57),
    .I1(1'b0),
    .I2(x37_y56),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001000110010)
) lut_40_61 (
    .O(x40_y61),
    .I0(x37_y62),
    .I1(x37_y61),
    .I2(x37_y57),
    .I3(x38_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011011110000)
) lut_41_61 (
    .O(x41_y61),
    .I0(x39_y62),
    .I1(1'b0),
    .I2(x39_y59),
    .I3(x39_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010101000010)
) lut_42_61 (
    .O(x42_y61),
    .I0(1'b0),
    .I1(x39_y57),
    .I2(x39_y62),
    .I3(x39_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101110111111)
) lut_43_61 (
    .O(x43_y61),
    .I0(x40_y61),
    .I1(x40_y57),
    .I2(x40_y62),
    .I3(x41_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001110011100)
) lut_44_61 (
    .O(x44_y61),
    .I0(1'b0),
    .I1(x42_y60),
    .I2(x42_y61),
    .I3(x42_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101011100111)
) lut_45_61 (
    .O(x45_y61),
    .I0(1'b0),
    .I1(x43_y61),
    .I2(x42_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011001100011)
) lut_46_61 (
    .O(x46_y61),
    .I0(x44_y60),
    .I1(x43_y59),
    .I2(x43_y62),
    .I3(x43_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111011001000)
) lut_47_61 (
    .O(x47_y61),
    .I0(1'b0),
    .I1(x45_y62),
    .I2(1'b0),
    .I3(x44_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010000100011)
) lut_48_61 (
    .O(x48_y61),
    .I0(x46_y61),
    .I1(x45_y59),
    .I2(x46_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110011000000)
) lut_49_61 (
    .O(x49_y61),
    .I0(x46_y60),
    .I1(1'b0),
    .I2(x47_y62),
    .I3(x46_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001010111000)
) lut_50_61 (
    .O(x50_y61),
    .I0(x48_y58),
    .I1(x48_y57),
    .I2(x48_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011101110001)
) lut_51_61 (
    .O(x51_y61),
    .I0(1'b0),
    .I1(x49_y62),
    .I2(1'b0),
    .I3(x49_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111101001011)
) lut_52_61 (
    .O(x52_y61),
    .I0(x50_y61),
    .I1(x49_y57),
    .I2(x50_y56),
    .I3(x50_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100000011001)
) lut_53_61 (
    .O(x53_y61),
    .I0(1'b0),
    .I1(x51_y59),
    .I2(x51_y59),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001000110011)
) lut_54_61 (
    .O(x54_y61),
    .I0(x51_y62),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x52_y56)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011010110001)
) lut_55_61 (
    .O(x55_y61),
    .I0(1'b0),
    .I1(x52_y62),
    .I2(x53_y61),
    .I3(x53_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001001111110)
) lut_56_61 (
    .O(x56_y61),
    .I0(x54_y58),
    .I1(x54_y62),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011010010110)
) lut_57_61 (
    .O(x57_y61),
    .I0(x55_y59),
    .I1(x55_y59),
    .I2(1'b0),
    .I3(x55_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110101101011)
) lut_58_61 (
    .O(x58_y61),
    .I0(x56_y62),
    .I1(1'b0),
    .I2(x56_y62),
    .I3(x56_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100011000000)
) lut_59_61 (
    .O(x59_y61),
    .I0(x56_y58),
    .I1(x56_y56),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111000011110)
) lut_60_61 (
    .O(x60_y61),
    .I0(1'b0),
    .I1(x58_y62),
    .I2(x58_y59),
    .I3(x58_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001100100101)
) lut_61_61 (
    .O(x61_y61),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x58_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010010000101)
) lut_62_61 (
    .O(x62_y61),
    .I0(1'b0),
    .I1(x59_y62),
    .I2(x59_y62),
    .I3(x60_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011010010111)
) lut_0_62 (
    .O(x0_y62),
    .I0(in2),
    .I1(in1),
    .I2(in2),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011011001110)
) lut_1_62 (
    .O(x1_y62),
    .I0(in2),
    .I1(in2),
    .I2(in2),
    .I3(in0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100110001101)
) lut_2_62 (
    .O(x2_y62),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001110001110)
) lut_3_62 (
    .O(x3_y62),
    .I0(in2),
    .I1(x1_y61),
    .I2(in1),
    .I3(x1_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011100101001)
) lut_4_62 (
    .O(x4_y62),
    .I0(1'b0),
    .I1(x1_y62),
    .I2(x2_y61),
    .I3(x1_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001100001100)
) lut_5_62 (
    .O(x5_y62),
    .I0(x2_y62),
    .I1(x2_y59),
    .I2(x3_y57),
    .I3(x2_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101100000110)
) lut_6_62 (
    .O(x6_y62),
    .I0(1'b0),
    .I1(x4_y62),
    .I2(x4_y57),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110111100010)
) lut_7_62 (
    .O(x7_y62),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x4_y62),
    .I3(x5_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011111001011)
) lut_8_62 (
    .O(x8_y62),
    .I0(x5_y62),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x5_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001100100001)
) lut_9_62 (
    .O(x9_y62),
    .I0(x6_y62),
    .I1(x6_y61),
    .I2(1'b0),
    .I3(x5_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000001111110)
) lut_10_62 (
    .O(x10_y62),
    .I0(1'b0),
    .I1(x7_y62),
    .I2(x7_y62),
    .I3(x8_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100011101001)
) lut_11_62 (
    .O(x11_y62),
    .I0(x9_y62),
    .I1(x8_y62),
    .I2(x8_y62),
    .I3(x9_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100111101101)
) lut_12_62 (
    .O(x12_y62),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x10_y62),
    .I3(x9_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001100101100)
) lut_13_62 (
    .O(x13_y62),
    .I0(x11_y62),
    .I1(x10_y60),
    .I2(x10_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111100001110)
) lut_14_62 (
    .O(x14_y62),
    .I0(x11_y62),
    .I1(x11_y62),
    .I2(x11_y62),
    .I3(x11_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011110111111)
) lut_15_62 (
    .O(x15_y62),
    .I0(x12_y61),
    .I1(x12_y61),
    .I2(x12_y60),
    .I3(x13_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010110111100)
) lut_16_62 (
    .O(x16_y62),
    .I0(x13_y61),
    .I1(1'b0),
    .I2(x14_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011110011100)
) lut_17_62 (
    .O(x17_y62),
    .I0(x14_y62),
    .I1(x15_y62),
    .I2(x15_y62),
    .I3(x14_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010111000101)
) lut_18_62 (
    .O(x18_y62),
    .I0(x16_y57),
    .I1(x16_y61),
    .I2(1'b0),
    .I3(x15_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101001101011)
) lut_19_62 (
    .O(x19_y62),
    .I0(x16_y62),
    .I1(x17_y59),
    .I2(x17_y61),
    .I3(x16_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101110001111)
) lut_20_62 (
    .O(x20_y62),
    .I0(x18_y61),
    .I1(x17_y62),
    .I2(1'b0),
    .I3(x18_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110011000000)
) lut_21_62 (
    .O(x21_y62),
    .I0(x19_y62),
    .I1(x18_y62),
    .I2(x18_y62),
    .I3(x19_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101110010110)
) lut_22_62 (
    .O(x22_y62),
    .I0(x20_y62),
    .I1(1'b0),
    .I2(x19_y61),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111000110100)
) lut_23_62 (
    .O(x23_y62),
    .I0(x21_y59),
    .I1(x20_y59),
    .I2(x21_y62),
    .I3(x21_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011100001111)
) lut_24_62 (
    .O(x24_y62),
    .I0(x21_y62),
    .I1(x22_y57),
    .I2(x21_y60),
    .I3(x21_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111011010100)
) lut_25_62 (
    .O(x25_y62),
    .I0(x23_y62),
    .I1(x22_y62),
    .I2(x23_y61),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010001000100)
) lut_26_62 (
    .O(x26_y62),
    .I0(x23_y62),
    .I1(x24_y60),
    .I2(x24_y58),
    .I3(x23_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101111001110)
) lut_27_62 (
    .O(x27_y62),
    .I0(x25_y62),
    .I1(x24_y59),
    .I2(x25_y61),
    .I3(x24_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000011110111)
) lut_28_62 (
    .O(x28_y62),
    .I0(1'b0),
    .I1(x25_y61),
    .I2(x26_y59),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010001101001)
) lut_29_62 (
    .O(x29_y62),
    .I0(x26_y62),
    .I1(x27_y62),
    .I2(x26_y58),
    .I3(x26_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010110100101)
) lut_30_62 (
    .O(x30_y62),
    .I0(x27_y62),
    .I1(x27_y62),
    .I2(x28_y57),
    .I3(x27_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111010001111)
) lut_31_62 (
    .O(x31_y62),
    .I0(1'b0),
    .I1(x29_y61),
    .I2(x28_y62),
    .I3(x29_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101101000011)
) lut_32_62 (
    .O(x32_y62),
    .I0(x30_y62),
    .I1(x29_y62),
    .I2(1'b0),
    .I3(x30_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111010110110)
) lut_33_62 (
    .O(x33_y62),
    .I0(1'b0),
    .I1(x30_y61),
    .I2(1'b0),
    .I3(x31_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110001111010)
) lut_34_62 (
    .O(x34_y62),
    .I0(x32_y58),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x32_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010101011110)
) lut_35_62 (
    .O(x35_y62),
    .I0(x33_y58),
    .I1(x32_y62),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010011100001)
) lut_36_62 (
    .O(x36_y62),
    .I0(x34_y60),
    .I1(x34_y58),
    .I2(1'b0),
    .I3(x33_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100110111010)
) lut_37_62 (
    .O(x37_y62),
    .I0(x34_y57),
    .I1(x35_y62),
    .I2(1'b0),
    .I3(x34_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111111011101)
) lut_38_62 (
    .O(x38_y62),
    .I0(1'b0),
    .I1(x35_y62),
    .I2(x36_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010110010000)
) lut_39_62 (
    .O(x39_y62),
    .I0(1'b0),
    .I1(x37_y59),
    .I2(x36_y57),
    .I3(x36_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111011011000)
) lut_40_62 (
    .O(x40_y62),
    .I0(x38_y62),
    .I1(1'b0),
    .I2(x37_y62),
    .I3(x38_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100011110111)
) lut_41_62 (
    .O(x41_y62),
    .I0(x39_y62),
    .I1(x38_y62),
    .I2(x39_y57),
    .I3(x38_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001101100100)
) lut_42_62 (
    .O(x42_y62),
    .I0(x39_y62),
    .I1(x39_y61),
    .I2(x39_y61),
    .I3(x40_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000100101001)
) lut_43_62 (
    .O(x43_y62),
    .I0(x40_y61),
    .I1(1'b0),
    .I2(x40_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010111100110)
) lut_44_62 (
    .O(x44_y62),
    .I0(x41_y62),
    .I1(x42_y62),
    .I2(x41_y58),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011010111011)
) lut_45_62 (
    .O(x45_y62),
    .I0(x42_y62),
    .I1(1'b0),
    .I2(x43_y62),
    .I3(x43_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011001000011)
) lut_46_62 (
    .O(x46_y62),
    .I0(x44_y62),
    .I1(x43_y62),
    .I2(x44_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011101100101)
) lut_47_62 (
    .O(x47_y62),
    .I0(x44_y62),
    .I1(1'b0),
    .I2(x44_y57),
    .I3(x44_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110101010000)
) lut_48_62 (
    .O(x48_y62),
    .I0(x45_y62),
    .I1(x46_y57),
    .I2(x46_y59),
    .I3(x46_y57)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110011100101)
) lut_49_62 (
    .O(x49_y62),
    .I0(x47_y57),
    .I1(x47_y62),
    .I2(x46_y60),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100101110011)
) lut_50_62 (
    .O(x50_y62),
    .I0(x47_y62),
    .I1(x47_y62),
    .I2(x47_y62),
    .I3(x47_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011100111000)
) lut_51_62 (
    .O(x51_y62),
    .I0(x48_y62),
    .I1(x48_y62),
    .I2(x49_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000110010010)
) lut_52_62 (
    .O(x52_y62),
    .I0(x50_y61),
    .I1(x49_y62),
    .I2(1'b0),
    .I3(x50_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111100010110)
) lut_53_62 (
    .O(x53_y62),
    .I0(x51_y62),
    .I1(x51_y62),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110011101111)
) lut_54_62 (
    .O(x54_y62),
    .I0(x52_y62),
    .I1(x52_y58),
    .I2(x52_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010000001110)
) lut_55_62 (
    .O(x55_y62),
    .I0(1'b0),
    .I1(x53_y62),
    .I2(x53_y62),
    .I3(x53_y61)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101100000101)
) lut_56_62 (
    .O(x56_y62),
    .I0(x54_y62),
    .I1(x53_y58),
    .I2(x53_y61),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000110110001)
) lut_57_62 (
    .O(x57_y62),
    .I0(x54_y62),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010000101111)
) lut_58_62 (
    .O(x58_y62),
    .I0(x56_y62),
    .I1(x55_y57),
    .I2(x55_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101001011101)
) lut_59_62 (
    .O(x59_y62),
    .I0(x57_y62),
    .I1(x57_y62),
    .I2(x57_y61),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001111011000)
) lut_60_62 (
    .O(x60_y62),
    .I0(1'b0),
    .I1(x57_y57),
    .I2(x58_y62),
    .I3(x57_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100011010111)
) lut_61_62 (
    .O(x61_y62),
    .I0(x58_y58),
    .I1(1'b0),
    .I2(x59_y58),
    .I3(x58_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111010010100)
) lut_62_62 (
    .O(x62_y62),
    .I0(x60_y59),
    .I1(1'b0),
    .I2(x60_y62),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000110101110)
) lut_0_63 (
    .O(x0_y63),
    .I0(in1),
    .I1(in2),
    .I2(1'b0),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100000000100)
) lut_1_63 (
    .O(x1_y63),
    .I0(in2),
    .I1(in1),
    .I2(in2),
    .I3(in1)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011001110101)
) lut_2_63 (
    .O(x2_y63),
    .I0(1'b0),
    .I1(in2),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010110111101)
) lut_3_63 (
    .O(x3_y63),
    .I0(x1_y61),
    .I1(1'b0),
    .I2(in1),
    .I3(in2)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110110101111)
) lut_4_63 (
    .O(x4_y63),
    .I0(x2_y62),
    .I1(x2_y61),
    .I2(x2_y58),
    .I3(x1_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011001111010)
) lut_5_63 (
    .O(x5_y63),
    .I0(x3_y61),
    .I1(x3_y62),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100000001110)
) lut_6_63 (
    .O(x6_y63),
    .I0(1'b0),
    .I1(x4_y62),
    .I2(1'b0),
    .I3(x4_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110011101011)
) lut_7_63 (
    .O(x7_y63),
    .I0(x5_y61),
    .I1(x5_y62),
    .I2(1'b0),
    .I3(x5_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111100100010)
) lut_8_63 (
    .O(x8_y63),
    .I0(x5_y62),
    .I1(x6_y62),
    .I2(x5_y62),
    .I3(x6_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110100111000)
) lut_9_63 (
    .O(x9_y63),
    .I0(x7_y62),
    .I1(x7_y58),
    .I2(x5_y62),
    .I3(x6_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011000001010)
) lut_10_63 (
    .O(x10_y63),
    .I0(1'b0),
    .I1(x8_y59),
    .I2(1'b0),
    .I3(x8_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010011000000)
) lut_11_63 (
    .O(x11_y63),
    .I0(1'b0),
    .I1(x8_y61),
    .I2(x8_y62),
    .I3(x9_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100000101011)
) lut_12_63 (
    .O(x12_y63),
    .I0(x10_y61),
    .I1(x9_y62),
    .I2(x10_y58),
    .I3(x9_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000110011010)
) lut_13_63 (
    .O(x13_y63),
    .I0(1'b0),
    .I1(x11_y59),
    .I2(x11_y61),
    .I3(x10_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100011000000)
) lut_14_63 (
    .O(x14_y63),
    .I0(x12_y62),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x11_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010101001001)
) lut_15_63 (
    .O(x15_y63),
    .I0(x12_y62),
    .I1(x12_y60),
    .I2(x12_y59),
    .I3(x12_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011111001111)
) lut_16_63 (
    .O(x16_y63),
    .I0(1'b0),
    .I1(x13_y62),
    .I2(x13_y60),
    .I3(1'b0)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011110100000)
) lut_17_63 (
    .O(x17_y63),
    .I0(x14_y59),
    .I1(1'b0),
    .I2(x14_y62),
    .I3(x15_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101110001110)
) lut_18_63 (
    .O(x18_y63),
    .I0(x15_y62),
    .I1(x15_y62),
    .I2(x16_y62),
    .I3(x15_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110011011111)
) lut_19_63 (
    .O(x19_y63),
    .I0(1'b0),
    .I1(x17_y62),
    .I2(x16_y62),
    .I3(x16_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011110001101)
) lut_20_63 (
    .O(x20_y63),
    .I0(x17_y62),
    .I1(x17_y60),
    .I2(x18_y62),
    .I3(x17_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100111000110)
) lut_21_63 (
    .O(x21_y63),
    .I0(x18_y62),
    .I1(x19_y62),
    .I2(1'b0),
    .I3(x19_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110011110101)
) lut_22_63 (
    .O(x22_y63),
    .I0(x19_y62),
    .I1(x20_y61),
    .I2(x19_y62),
    .I3(x20_y60)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011010001100)
) lut_23_63 (
    .O(x23_y63),
    .I0(x21_y62),
    .I1(x20_y62),
    .I2(1'b0),
    .I3(x20_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101111100101)
) lut_24_63 (
    .O(x24_y63),
    .I0(x22_y62),
    .I1(x22_y61),
    .I2(x21_y60),
    .I3(x22_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100101001011)
) lut_25_63 (
    .O(x25_y63),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x22_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011000111010)
) lut_26_63 (
    .O(x26_y63),
    .I0(x24_y62),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x24_y58)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011001110010)
) lut_27_63 (
    .O(x27_y63),
    .I0(x25_y59),
    .I1(1'b0),
    .I2(x24_y62),
    .I3(x25_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001101011000)
) lut_28_63 (
    .O(x28_y63),
    .I0(x25_y62),
    .I1(x25_y62),
    .I2(x26_y58),
    .I3(x26_y62)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010100111011)
) lut_29_63 (
    .O(x29_y63),
    .I0(x27_y62),
    .I1(x26_y62),
    .I2(x26_y62),
    .I3(x27_y59)
);

(* keep, dont_touch *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010100010001)
) lut_30_63 (
    .O(x30_y63),
    .I0(x27_y62),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

endmodule