module individual (
    (* keep *) input in0, in1, in2, in3, in4, in5, in6, in7, in8, in9,
    (* keep *) output out0, out1, out2, out3, out4, out5, out6, out7, out8, out9);
    wire x1_y1;
    wire x2_y1;
    wire x3_y1;
    wire x4_y1;
    wire x5_y1;
    wire x7_y1;
    wire x8_y1;
    wire x9_y1;
    wire x10_y1;
    wire x11_y1;
    wire x1_y2;
    wire x2_y2;
    wire x3_y2;
    wire x4_y2;
    wire x5_y2;
    wire x7_y2;
    wire x8_y2;
    wire x9_y2;
    wire x10_y2;
    wire x11_y2;
    wire x1_y3;
    wire x2_y3;
    wire x3_y3;
    wire x4_y3;
    wire x5_y3;
    wire x7_y3;
    wire x8_y3;
    wire x9_y3;
    wire x10_y3;
    wire x11_y3;
    wire x1_y4;
    wire x2_y4;
    wire x3_y4;
    wire x4_y4;
    wire x5_y4;
    wire x7_y4;
    wire x8_y4;
    wire x9_y4;
    wire x10_y4;
    wire x11_y4;
    wire x1_y5;
    wire x2_y5;
    wire x3_y5;
    wire x4_y5;
    wire x5_y5;
    wire x7_y5;
    wire x8_y5;
    wire x9_y5;
    wire x10_y5;
    wire x11_y5;
    wire x1_y6;
    wire x2_y6;
    wire x3_y6;
    wire x4_y6;
    wire x5_y6;
    wire x7_y6;
    wire x8_y6;
    wire x9_y6;
    wire x10_y6;
    wire x11_y6;
    wire x1_y7;
    wire x2_y7;
    wire x3_y7;
    wire x4_y7;
    wire x5_y7;
    wire x7_y7;
    wire x8_y7;
    wire x9_y7;
    wire x10_y7;
    wire x11_y7;
    wire x1_y8;
    wire x2_y8;
    wire x3_y8;
    wire x4_y8;
    wire x5_y8;
    wire x7_y8;
    wire x8_y8;
    wire x9_y8;
    wire x10_y8;
    wire x11_y8;
    wire x1_y9;
    wire x2_y9;
    wire x3_y9;
    wire x4_y9;
    wire x5_y9;
    wire x7_y9;
    wire x8_y9;
    wire x9_y9;
    wire x10_y9;
    wire x11_y9;
    wire x1_y10;
    wire x2_y10;
    wire x3_y10;
    wire x4_y10;
    wire x5_y10;
    wire x7_y10;
    wire x8_y10;
    wire x9_y10;
    wire x10_y10;
    wire x11_y10;

    (* keep, dont_touch *)
    (* BEL = "X1/Y1/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000111)
    ) lut_0 (
        .O(out_0),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X2/Y1/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001000)
    ) lut_1 (
        .O(out_1),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X3/Y1/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001000)
    ) lut_2 (
        .O(out_2),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X4/Y1/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000111)
    ) lut_3 (
        .O(out_3),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X5/Y1/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001111)
    ) lut_4 (
        .O(out_4),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X7/Y1/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000101)
    ) lut_5 (
        .O(out_5),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X8/Y1/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001001)
    ) lut_6 (
        .O(out_6),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X9/Y1/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000001)
    ) lut_7 (
        .O(out_7),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X10/Y1/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001111)
    ) lut_8 (
        .O(out_8),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X11/Y1/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000001)
    ) lut_9 (
        .O(out_9),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X1/Y1/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001001)
    ) lut_10 (
        .O(out_10),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X2/Y1/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000010)
    ) lut_11 (
        .O(out_11),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X3/Y1/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001010)
    ) lut_12 (
        .O(out_12),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X4/Y1/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000101)
    ) lut_13 (
        .O(out_13),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X5/Y1/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001010)
    ) lut_14 (
        .O(out_14),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X7/Y1/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000110)
    ) lut_15 (
        .O(out_15),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X8/Y1/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000011)
    ) lut_16 (
        .O(out_16),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X9/Y1/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000011)
    ) lut_17 (
        .O(out_17),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X10/Y1/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001100)
    ) lut_18 (
        .O(out_18),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X11/Y1/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001110)
    ) lut_19 (
        .O(out_19),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X1/Y1/lc2" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001101)
    ) lut_20 (
        .O(out_20),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X2/Y1/lc2" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001110)
    ) lut_21 (
        .O(out_21),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X3/Y1/lc2" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001001)
    ) lut_22 (
        .O(out_22),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X4/Y1/lc2" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001010)
    ) lut_23 (
        .O(out_23),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X5/Y1/lc2" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000100)
    ) lut_24 (
        .O(out_24),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X7/Y1/lc2" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000000)
    ) lut_25 (
        .O(out_25),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X8/Y1/lc2" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000110)
    ) lut_26 (
        .O(out_26),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X9/Y1/lc2" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001101)
    ) lut_27 (
        .O(out_27),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X10/Y1/lc2" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001110)
    ) lut_28 (
        .O(out_28),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X11/Y1/lc2" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001110)
    ) lut_29 (
        .O(out_29),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X1/Y1/lc3" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000100)
    ) lut_30 (
        .O(out_30),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X2/Y1/lc3" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000111)
    ) lut_31 (
        .O(out_31),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X3/Y1/lc3" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001011)
    ) lut_32 (
        .O(out_32),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X4/Y1/lc3" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000110)
    ) lut_33 (
        .O(out_33),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X5/Y1/lc3" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001010)
    ) lut_34 (
        .O(out_34),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X7/Y1/lc3" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000110)
    ) lut_35 (
        .O(out_35),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X8/Y1/lc3" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001001)
    ) lut_36 (
        .O(out_36),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X9/Y1/lc3" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000001)
    ) lut_37 (
        .O(out_37),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X10/Y1/lc3" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000000)
    ) lut_38 (
        .O(out_38),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X11/Y1/lc3" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001110)
    ) lut_39 (
        .O(out_39),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X1/Y1/lc4" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001100)
    ) lut_40 (
        .O(out_40),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X2/Y1/lc4" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000111)
    ) lut_41 (
        .O(out_41),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X3/Y1/lc4" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000001)
    ) lut_42 (
        .O(out_42),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X4/Y1/lc4" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000011)
    ) lut_43 (
        .O(out_43),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X5/Y1/lc4" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000111)
    ) lut_44 (
        .O(out_44),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X7/Y1/lc4" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001111)
    ) lut_45 (
        .O(out_45),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X8/Y1/lc4" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001000)
    ) lut_46 (
        .O(out_46),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X9/Y1/lc4" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001101)
    ) lut_47 (
        .O(out_47),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X10/Y1/lc4" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000000)
    ) lut_48 (
        .O(out_48),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X11/Y1/lc4" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001110)
    ) lut_49 (
        .O(out_49),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X1/Y1/lc5" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000100)
    ) lut_50 (
        .O(out_50),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X2/Y1/lc5" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000001)
    ) lut_51 (
        .O(out_51),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X3/Y1/lc5" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001011)
    ) lut_52 (
        .O(out_52),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X4/Y1/lc5" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000111)
    ) lut_53 (
        .O(out_53),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X5/Y1/lc5" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000101)
    ) lut_54 (
        .O(out_54),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X7/Y1/lc5" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000101)
    ) lut_55 (
        .O(out_55),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X8/Y1/lc5" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001000)
    ) lut_56 (
        .O(out_56),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X9/Y1/lc5" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001101)
    ) lut_57 (
        .O(out_57),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X10/Y1/lc5" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000001)
    ) lut_58 (
        .O(out_58),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X11/Y1/lc5" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001111)
    ) lut_59 (
        .O(out_59),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X1/Y1/lc6" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000101)
    ) lut_60 (
        .O(out_60),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X2/Y1/lc6" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001100)
    ) lut_61 (
        .O(out_61),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X3/Y1/lc6" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001011)
    ) lut_62 (
        .O(out_62),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X4/Y1/lc6" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001010)
    ) lut_63 (
        .O(out_63),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X5/Y1/lc6" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000011)
    ) lut_64 (
        .O(out_64),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X7/Y1/lc6" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001010)
    ) lut_65 (
        .O(out_65),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X8/Y1/lc6" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001101)
    ) lut_66 (
        .O(out_66),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X9/Y1/lc6" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000000)
    ) lut_67 (
        .O(out_67),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X10/Y1/lc6" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001000)
    ) lut_68 (
        .O(out_68),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X11/Y1/lc6" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000110)
    ) lut_69 (
        .O(out_69),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X1/Y1/lc7" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001001)
    ) lut_70 (
        .O(out_70),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X2/Y1/lc7" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000010)
    ) lut_71 (
        .O(out_71),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X3/Y1/lc7" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000011)
    ) lut_72 (
        .O(out_72),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X4/Y1/lc7" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000111)
    ) lut_73 (
        .O(out_73),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X5/Y1/lc7" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001001)
    ) lut_74 (
        .O(out_74),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X7/Y1/lc7" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000011)
    ) lut_75 (
        .O(out_75),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X8/Y1/lc7" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001101)
    ) lut_76 (
        .O(out_76),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X9/Y1/lc7" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001111)
    ) lut_77 (
        .O(out_77),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X10/Y1/lc7" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000101)
    ) lut_78 (
        .O(out_78),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X11/Y1/lc7" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001110)
    ) lut_79 (
        .O(out_79),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X1/Y2/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001101)
    ) lut_80 (
        .O(out_80),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X2/Y2/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000111)
    ) lut_81 (
        .O(out_81),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X3/Y2/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000010)
    ) lut_82 (
        .O(out_82),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X4/Y2/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001011)
    ) lut_83 (
        .O(out_83),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X5/Y2/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000100)
    ) lut_84 (
        .O(out_84),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X7/Y2/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001000)
    ) lut_85 (
        .O(out_85),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X8/Y2/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001111)
    ) lut_86 (
        .O(out_86),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X9/Y2/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001010)
    ) lut_87 (
        .O(out_87),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X10/Y2/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001100)
    ) lut_88 (
        .O(out_88),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X11/Y2/lc0" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001110)
    ) lut_89 (
        .O(out_89),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X1/Y2/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001010)
    ) lut_90 (
        .O(out_90),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X2/Y2/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001101)
    ) lut_91 (
        .O(out_91),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X3/Y2/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001011)
    ) lut_92 (
        .O(out_92),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X4/Y2/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000111)
    ) lut_93 (
        .O(out_93),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X5/Y2/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000001)
    ) lut_94 (
        .O(out_94),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X7/Y2/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000110)
    ) lut_95 (
        .O(out_95),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X8/Y2/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000111)
    ) lut_96 (
        .O(out_96),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X9/Y2/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001101)
    ) lut_97 (
        .O(out_97),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X10/Y2/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000001010)
    ) lut_98 (
        .O(out_98),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
    (* keep, dont_touch *)
    (* BEL = "X11/Y2/lc1" *)
    SB_LUT4 #(
        .LUT_INIT(16'b0000000000000011)
    ) lut_99 (
        .O(out_99),
        .I0(/* input0 connection */),
        .I1(/* input1 connection */),
        .I2(/* input2 connection */),
        .I3(/* input3 connection */)
    );
endmodule
