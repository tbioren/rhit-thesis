module cgp_module (
    (* keep *) input in0, in1, in2, in3, in4, in5, in6, in7, in8, in9,
    (* keep *) output out0, out1, out2, out3, out4, out5, out6, out7, out8, out9);

    (* keep *) wire x0_y0, x1_y0, x2_y0, x3_y0, x4_y0, x5_y0, x6_y0, x7_y0, x8_y0, x9_y0, x10_y0, x11_y0, x12_y0, x13_y0, x14_y0, x15_y0, x16_y0, x17_y0, x18_y0, x19_y0, x20_y0, x21_y0, x22_y0, x23_y0, x24_y0, x25_y0, x26_y0, x27_y0, x28_y0, x29_y0, x30_y0, x31_y0, x32_y0, x33_y0, x34_y0, x35_y0, x36_y0, x37_y0, x38_y0, x39_y0, x40_y0, x41_y0, x42_y0, x43_y0, x44_y0, x45_y0, x46_y0, x47_y0, x48_y0, x0_y1, x1_y1, x2_y1, x3_y1, x4_y1, x5_y1, x6_y1, x7_y1, x8_y1, x9_y1, x10_y1, x11_y1, x12_y1, x13_y1, x14_y1, x15_y1, x16_y1, x17_y1, x18_y1, x19_y1, x20_y1, x21_y1, x22_y1, x23_y1, x24_y1, x25_y1, x26_y1, x27_y1, x28_y1, x29_y1, x30_y1, x31_y1, x32_y1, x33_y1, x34_y1, x35_y1, x36_y1, x37_y1, x38_y1, x39_y1, x40_y1, x41_y1, x42_y1, x43_y1, x44_y1, x45_y1, x46_y1, x47_y1, x48_y1, x0_y2, x1_y2, x2_y2, x3_y2, x4_y2, x5_y2, x6_y2, x7_y2, x8_y2, x9_y2, x10_y2, x11_y2, x12_y2, x13_y2, x14_y2, x15_y2, x16_y2, x17_y2, x18_y2, x19_y2, x20_y2, x21_y2, x22_y2, x23_y2, x24_y2, x25_y2, x26_y2, x27_y2, x28_y2, x29_y2, x30_y2, x31_y2, x32_y2, x33_y2, x34_y2, x35_y2, x36_y2, x37_y2, x38_y2, x39_y2, x40_y2, x41_y2, x42_y2, x43_y2, x44_y2, x45_y2, x46_y2, x47_y2, x48_y2, x0_y3, x1_y3, x2_y3, x3_y3, x4_y3, x5_y3, x6_y3, x7_y3, x8_y3, x9_y3, x10_y3, x11_y3, x12_y3, x13_y3, x14_y3, x15_y3, x16_y3, x17_y3, x18_y3, x19_y3, x20_y3, x21_y3, x22_y3, x23_y3, x24_y3, x25_y3, x26_y3, x27_y3, x28_y3, x29_y3, x30_y3, x31_y3, x32_y3, x33_y3, x34_y3, x35_y3, x36_y3, x37_y3, x38_y3, x39_y3, x40_y3, x41_y3, x42_y3, x43_y3, x44_y3, x45_y3, x46_y3, x47_y3, x48_y3, x0_y4, x1_y4, x2_y4, x3_y4, x4_y4, x5_y4, x6_y4, x7_y4, x8_y4, x9_y4, x10_y4, x11_y4, x12_y4, x13_y4, x14_y4, x15_y4, x16_y4, x17_y4, x18_y4, x19_y4, x20_y4, x21_y4, x22_y4, x23_y4, x24_y4, x25_y4, x26_y4, x27_y4, x28_y4, x29_y4, x30_y4, x31_y4, x32_y4, x33_y4, x34_y4, x35_y4, x36_y4, x37_y4, x38_y4, x39_y4, x40_y4, x41_y4, x42_y4, x43_y4, x44_y4, x45_y4, x46_y4, x47_y4, x48_y4, x0_y5, x1_y5, x2_y5, x3_y5, x4_y5, x5_y5, x6_y5, x7_y5, x8_y5, x9_y5, x10_y5, x11_y5, x12_y5, x13_y5, x14_y5, x15_y5, x16_y5, x17_y5, x18_y5, x19_y5, x20_y5, x21_y5, x22_y5, x23_y5, x24_y5, x25_y5, x26_y5, x27_y5, x28_y5, x29_y5, x30_y5, x31_y5, x32_y5, x33_y5, x34_y5, x35_y5, x36_y5, x37_y5, x38_y5, x39_y5, x40_y5, x41_y5, x42_y5, x43_y5, x44_y5, x45_y5, x46_y5, x47_y5, x48_y5, x0_y6, x1_y6, x2_y6, x3_y6, x4_y6, x5_y6, x6_y6, x7_y6, x8_y6, x9_y6, x10_y6, x11_y6, x12_y6, x13_y6, x14_y6, x15_y6, x16_y6, x17_y6, x18_y6, x19_y6, x20_y6, x21_y6, x22_y6, x23_y6, x24_y6, x25_y6, x26_y6, x27_y6, x28_y6, x29_y6, x30_y6, x31_y6, x32_y6, x33_y6, x34_y6, x35_y6, x36_y6, x37_y6, x38_y6, x39_y6, x40_y6, x41_y6, x42_y6, x43_y6, x44_y6, x45_y6, x46_y6, x47_y6, x48_y6, x0_y7, x1_y7, x2_y7, x3_y7, x4_y7, x5_y7, x6_y7, x7_y7, x8_y7, x9_y7, x10_y7, x11_y7, x12_y7, x13_y7, x14_y7, x15_y7, x16_y7, x17_y7, x18_y7, x19_y7, x20_y7, x21_y7, x22_y7, x23_y7, x24_y7, x25_y7, x26_y7, x27_y7, x28_y7, x29_y7, x30_y7, x31_y7, x32_y7, x33_y7, x34_y7, x35_y7, x36_y7, x37_y7, x38_y7, x39_y7, x40_y7, x41_y7, x42_y7, x43_y7, x44_y7, x45_y7, x46_y7, x47_y7, x48_y7, x0_y8, x1_y8, x2_y8, x3_y8, x4_y8, x5_y8, x6_y8, x7_y8, x8_y8, x9_y8, x10_y8, x11_y8, x12_y8, x13_y8, x14_y8, x15_y8, x16_y8, x17_y8, x18_y8, x19_y8, x20_y8, x21_y8, x22_y8, x23_y8, x24_y8, x25_y8, x26_y8, x27_y8, x28_y8, x29_y8, x30_y8, x31_y8, x32_y8, x33_y8, x34_y8, x35_y8, x36_y8, x37_y8, x38_y8, x39_y8, x40_y8, x41_y8, x42_y8, x43_y8, x44_y8, x45_y8, x46_y8, x47_y8, x48_y8, x0_y9, x1_y9, x2_y9, x3_y9, x4_y9, x5_y9, x6_y9, x7_y9, x8_y9, x9_y9, x10_y9, x11_y9, x12_y9, x13_y9, x14_y9, x15_y9, x16_y9, x17_y9, x18_y9, x19_y9, x20_y9, x21_y9, x22_y9, x23_y9, x24_y9, x25_y9, x26_y9, x27_y9, x28_y9, x29_y9, x30_y9, x31_y9, x32_y9, x33_y9, x34_y9, x35_y9, x36_y9, x37_y9, x38_y9, x39_y9, x40_y9, x41_y9, x42_y9, x43_y9, x44_y9, x45_y9, x46_y9, x47_y9, x48_y9, x0_y10, x1_y10, x2_y10, x3_y10, x4_y10, x5_y10, x6_y10, x7_y10, x8_y10, x9_y10, x10_y10, x11_y10, x12_y10, x13_y10, x14_y10, x15_y10, x16_y10, x17_y10, x18_y10, x19_y10, x20_y10, x21_y10, x22_y10, x23_y10, x24_y10, x25_y10, x26_y10, x27_y10, x28_y10, x29_y10, x30_y10, x31_y10, x32_y10, x33_y10, x34_y10, x35_y10, x36_y10, x37_y10, x38_y10, x39_y10, x40_y10, x41_y10, x42_y10, x43_y10, x44_y10, x45_y10, x46_y10, x47_y10, x48_y10, x0_y11, x1_y11, x2_y11, x3_y11, x4_y11, x5_y11, x6_y11, x7_y11, x8_y11, x9_y11, x10_y11, x11_y11, x12_y11, x13_y11, x14_y11, x15_y11, x16_y11, x17_y11, x18_y11, x19_y11, x20_y11, x21_y11, x22_y11, x23_y11, x24_y11, x25_y11, x26_y11, x27_y11, x28_y11, x29_y11, x30_y11, x31_y11, x32_y11, x33_y11, x34_y11, x35_y11, x36_y11, x37_y11, x38_y11, x39_y11, x40_y11, x41_y11, x42_y11, x43_y11, x44_y11, x45_y11, x46_y11, x47_y11, x48_y11, x0_y12, x1_y12, x2_y12, x3_y12, x4_y12, x5_y12, x6_y12, x7_y12, x8_y12, x9_y12, x10_y12, x11_y12, x12_y12, x13_y12, x14_y12, x15_y12, x16_y12, x17_y12, x18_y12, x19_y12, x20_y12, x21_y12, x22_y12, x23_y12, x24_y12, x25_y12, x26_y12, x27_y12, x28_y12, x29_y12, x30_y12, x31_y12, x32_y12, x33_y12, x34_y12, x35_y12, x36_y12, x37_y12, x38_y12, x39_y12, x40_y12, x41_y12, x42_y12, x43_y12, x44_y12, x45_y12, x46_y12, x47_y12, x48_y12, x0_y13, x1_y13, x2_y13, x3_y13, x4_y13, x5_y13, x6_y13, x7_y13, x8_y13, x9_y13, x10_y13, x11_y13, x12_y13, x13_y13, x14_y13, x15_y13, x16_y13, x17_y13, x18_y13, x19_y13, x20_y13, x21_y13, x22_y13, x23_y13, x24_y13, x25_y13, x26_y13, x27_y13, x28_y13, x29_y13, x30_y13, x31_y13, x32_y13, x33_y13, x34_y13, x35_y13, x36_y13, x37_y13, x38_y13, x39_y13, x40_y13, x41_y13, x42_y13, x43_y13, x44_y13, x45_y13, x46_y13, x47_y13, x48_y13, x0_y14, x1_y14, x2_y14, x3_y14, x4_y14, x5_y14, x6_y14, x7_y14, x8_y14, x9_y14, x10_y14, x11_y14, x12_y14, x13_y14, x14_y14, x15_y14, x16_y14, x17_y14, x18_y14, x19_y14, x20_y14, x21_y14, x22_y14, x23_y14, x24_y14, x25_y14, x26_y14, x27_y14, x28_y14, x29_y14, x30_y14, x31_y14, x32_y14, x33_y14, x34_y14, x35_y14, x36_y14, x37_y14, x38_y14, x39_y14, x40_y14, x41_y14, x42_y14, x43_y14, x44_y14, x45_y14, x46_y14, x47_y14, x48_y14, x0_y15, x1_y15, x2_y15, x3_y15, x4_y15, x5_y15, x6_y15, x7_y15, x8_y15, x9_y15, x10_y15, x11_y15, x12_y15, x13_y15, x14_y15, x15_y15, x16_y15, x17_y15, x18_y15, x19_y15, x20_y15, x21_y15, x22_y15, x23_y15, x24_y15, x25_y15, x26_y15, x27_y15, x28_y15, x29_y15, x30_y15, x31_y15, x32_y15, x33_y15, x34_y15, x35_y15, x36_y15, x37_y15, x38_y15, x39_y15, x40_y15, x41_y15, x42_y15, x43_y15, x44_y15, x45_y15, x46_y15, x47_y15, x48_y15, x0_y16, x1_y16, x2_y16, x3_y16, x4_y16, x5_y16, x6_y16, x7_y16, x8_y16, x9_y16, x10_y16, x11_y16, x12_y16, x13_y16, x14_y16, x15_y16, x16_y16, x17_y16, x18_y16, x19_y16, x20_y16, x21_y16, x22_y16, x23_y16, x24_y16, x25_y16, x26_y16, x27_y16, x28_y16, x29_y16, x30_y16, x31_y16, x32_y16, x33_y16, x34_y16, x35_y16, x36_y16, x37_y16, x38_y16, x39_y16, x40_y16, x41_y16, x42_y16, x43_y16, x44_y16, x45_y16, x46_y16, x47_y16, x48_y16, x0_y17, x1_y17, x2_y17, x3_y17, x4_y17, x5_y17, x6_y17, x7_y17, x8_y17, x9_y17, x10_y17, x11_y17, x12_y17, x13_y17, x14_y17, x15_y17, x16_y17, x17_y17, x18_y17, x19_y17, x20_y17, x21_y17, x22_y17, x23_y17, x24_y17, x25_y17, x26_y17, x27_y17, x28_y17, x29_y17, x30_y17, x31_y17, x32_y17, x33_y17, x34_y17, x35_y17, x36_y17, x37_y17, x38_y17, x39_y17, x40_y17, x41_y17, x42_y17, x43_y17, x44_y17, x45_y17, x46_y17, x47_y17, x48_y17, x0_y18, x1_y18, x2_y18, x3_y18, x4_y18, x5_y18, x6_y18, x7_y18, x8_y18, x9_y18, x10_y18, x11_y18, x12_y18, x13_y18, x14_y18, x15_y18, x16_y18, x17_y18, x18_y18, x19_y18, x20_y18, x21_y18, x22_y18, x23_y18, x24_y18, x25_y18, x26_y18, x27_y18, x28_y18, x29_y18, x30_y18, x31_y18, x32_y18, x33_y18, x34_y18, x35_y18, x36_y18, x37_y18, x38_y18, x39_y18, x40_y18, x41_y18, x42_y18, x43_y18, x44_y18, x45_y18, x46_y18, x47_y18, x48_y18, x0_y19, x1_y19, x2_y19, x3_y19, x4_y19, x5_y19, x6_y19, x7_y19, x8_y19, x9_y19, x10_y19, x11_y19, x12_y19, x13_y19, x14_y19, x15_y19, x16_y19, x17_y19, x18_y19, x19_y19, x20_y19, x21_y19, x22_y19, x23_y19, x24_y19, x25_y19, x26_y19, x27_y19, x28_y19, x29_y19, x30_y19, x31_y19, x32_y19, x33_y19, x34_y19, x35_y19, x36_y19, x37_y19, x38_y19, x39_y19, x40_y19, x41_y19, x42_y19, x43_y19, x44_y19, x45_y19, x46_y19, x47_y19, x48_y19, x0_y20, x1_y20, x2_y20, x3_y20, x4_y20, x5_y20, x6_y20, x7_y20, x8_y20, x9_y20, x10_y20, x11_y20, x12_y20, x13_y20, x14_y20, x15_y20, x16_y20, x17_y20, x18_y20, x19_y20, x20_y20, x21_y20, x22_y20, x23_y20, x24_y20, x25_y20, x26_y20, x27_y20, x28_y20, x29_y20, x30_y20, x31_y20, x32_y20, x33_y20, x34_y20, x35_y20, x36_y20, x37_y20, x38_y20, x39_y20, x40_y20, x41_y20, x42_y20, x43_y20, x44_y20, x45_y20, x46_y20, x47_y20, x48_y20, x0_y21, x1_y21, x2_y21, x3_y21, x4_y21, x5_y21, x6_y21, x7_y21, x8_y21, x9_y21, x10_y21, x11_y21, x12_y21, x13_y21, x14_y21, x15_y21, x16_y21, x17_y21, x18_y21, x19_y21, x20_y21, x21_y21, x22_y21, x23_y21, x24_y21, x25_y21, x26_y21, x27_y21, x28_y21, x29_y21, x30_y21, x31_y21, x32_y21, x33_y21, x34_y21, x35_y21, x36_y21, x37_y21, x38_y21, x39_y21, x40_y21, x41_y21, x42_y21, x43_y21, x44_y21, x45_y21, x46_y21, x47_y21, x48_y21, x0_y22, x1_y22, x2_y22, x3_y22, x4_y22, x5_y22, x6_y22, x7_y22, x8_y22, x9_y22, x10_y22, x11_y22, x12_y22, x13_y22, x14_y22, x15_y22, x16_y22, x17_y22, x18_y22, x19_y22, x20_y22, x21_y22, x22_y22, x23_y22, x24_y22, x25_y22, x26_y22, x27_y22, x28_y22, x29_y22, x30_y22, x31_y22, x32_y22, x33_y22, x34_y22, x35_y22, x36_y22, x37_y22, x38_y22, x39_y22, x40_y22, x41_y22, x42_y22, x43_y22, x44_y22, x45_y22, x46_y22, x47_y22, x48_y22, x0_y23, x1_y23, x2_y23, x3_y23, x4_y23, x5_y23, x6_y23, x7_y23, x8_y23, x9_y23, x10_y23, x11_y23, x12_y23, x13_y23, x14_y23, x15_y23, x16_y23, x17_y23, x18_y23, x19_y23, x20_y23, x21_y23, x22_y23, x23_y23, x24_y23, x25_y23, x26_y23, x27_y23, x28_y23, x29_y23, x30_y23, x31_y23, x32_y23, x33_y23, x34_y23, x35_y23, x36_y23, x37_y23, x38_y23, x39_y23, x40_y23, x41_y23, x42_y23, x43_y23, x44_y23, x45_y23, x46_y23, x47_y23, x48_y23, x0_y24, x1_y24, x2_y24, x3_y24, x4_y24, x5_y24, x6_y24, x7_y24, x8_y24, x9_y24, x10_y24, x11_y24, x12_y24, x13_y24, x14_y24, x15_y24, x16_y24, x17_y24, x18_y24, x19_y24, x20_y24, x21_y24, x22_y24, x23_y24, x24_y24, x25_y24, x26_y24, x27_y24, x28_y24, x29_y24, x30_y24, x31_y24, x32_y24, x33_y24, x34_y24, x35_y24, x36_y24, x37_y24, x38_y24, x39_y24, x40_y24, x41_y24, x42_y24, x43_y24, x44_y24, x45_y24, x46_y24, x47_y24, x48_y24, x0_y25, x1_y25, x2_y25, x3_y25, x4_y25, x5_y25, x6_y25, x7_y25, x8_y25, x9_y25, x10_y25, x11_y25, x12_y25, x13_y25, x14_y25, x15_y25, x16_y25, x17_y25, x18_y25, x19_y25, x20_y25, x21_y25, x22_y25, x23_y25, x24_y25, x25_y25, x26_y25, x27_y25, x28_y25, x29_y25, x30_y25, x31_y25, x32_y25, x33_y25, x34_y25, x35_y25, x36_y25, x37_y25, x38_y25, x39_y25, x40_y25, x41_y25, x42_y25, x43_y25, x44_y25, x45_y25, x46_y25, x47_y25, x48_y25, x0_y26, x1_y26, x2_y26, x3_y26, x4_y26, x5_y26, x6_y26, x7_y26, x8_y26, x9_y26, x10_y26, x11_y26, x12_y26, x13_y26, x14_y26, x15_y26, x16_y26, x17_y26, x18_y26, x19_y26, x20_y26, x21_y26, x22_y26, x23_y26, x24_y26, x25_y26, x26_y26, x27_y26, x28_y26, x29_y26, x30_y26, x31_y26, x32_y26, x33_y26, x34_y26, x35_y26, x36_y26, x37_y26, x38_y26, x39_y26, x40_y26, x41_y26, x42_y26, x43_y26, x44_y26, x45_y26, x46_y26, x47_y26, x48_y26, x0_y27, x1_y27, x2_y27, x3_y27, x4_y27, x5_y27, x6_y27, x7_y27, x8_y27, x9_y27, x10_y27, x11_y27, x12_y27, x13_y27, x14_y27, x15_y27, x16_y27, x17_y27, x18_y27, x19_y27, x20_y27, x21_y27, x22_y27, x23_y27, x24_y27, x25_y27, x26_y27, x27_y27, x28_y27, x29_y27, x30_y27, x31_y27, x32_y27, x33_y27, x34_y27, x35_y27, x36_y27, x37_y27, x38_y27, x39_y27, x40_y27, x41_y27, x42_y27, x43_y27, x44_y27, x45_y27, x46_y27, x47_y27, x48_y27, x0_y28, x1_y28, x2_y28, x3_y28, x4_y28, x5_y28, x6_y28, x7_y28, x8_y28, x9_y28, x10_y28, x11_y28, x12_y28, x13_y28, x14_y28, x15_y28, x16_y28, x17_y28, x18_y28, x19_y28, x20_y28, x21_y28, x22_y28, x23_y28, x24_y28, x25_y28, x26_y28, x27_y28, x28_y28, x29_y28, x30_y28, x31_y28, x32_y28, x33_y28, x34_y28, x35_y28, x36_y28, x37_y28, x38_y28, x39_y28, x40_y28, x41_y28, x42_y28, x43_y28, x44_y28, x45_y28, x46_y28, x47_y28, x48_y28, x0_y29, x1_y29, x2_y29, x3_y29, x4_y29, x5_y29, x6_y29, x7_y29, x8_y29, x9_y29, x10_y29, x11_y29, x12_y29, x13_y29, x14_y29, x15_y29, x16_y29, x17_y29, x18_y29, x19_y29, x20_y29, x21_y29, x22_y29, x23_y29, x24_y29, x25_y29, x26_y29, x27_y29, x28_y29, x29_y29, x30_y29, x31_y29, x32_y29, x33_y29, x34_y29, x35_y29, x36_y29, x37_y29, x38_y29, x39_y29, x40_y29, x41_y29, x42_y29, x43_y29, x44_y29, x45_y29, x46_y29, x47_y29, x48_y29, x0_y30, x1_y30, x2_y30, x3_y30, x4_y30, x5_y30, x6_y30, x7_y30, x8_y30, x9_y30, x10_y30, x11_y30, x12_y30, x13_y30, x14_y30, x15_y30, x16_y30, x17_y30, x18_y30, x19_y30, x20_y30, x21_y30, x22_y30, x23_y30, x24_y30, x25_y30, x26_y30, x27_y30, x28_y30, x29_y30, x30_y30, x31_y30, x32_y30, x33_y30, x34_y30, x35_y30, x36_y30, x37_y30, x38_y30, x39_y30, x40_y30, x41_y30, x42_y30, x43_y30, x44_y30, x45_y30, x46_y30, x47_y30, x48_y30, x0_y31, x1_y31, x2_y31, x3_y31, x4_y31, x5_y31, x6_y31, x7_y31, x8_y31, x9_y31, x10_y31, x11_y31, x12_y31, x13_y31, x14_y31, x15_y31, x16_y31, x17_y31, x18_y31, x19_y31, x20_y31, x21_y31, x22_y31, x23_y31, x24_y31, x25_y31, x26_y31, x27_y31, x28_y31, x29_y31, x30_y31, x31_y31, x32_y31, x33_y31, x34_y31, x35_y31, x36_y31, x37_y31, x38_y31, x39_y31, x40_y31, x41_y31, x42_y31, x43_y31, x44_y31, x45_y31, x46_y31, x47_y31, x48_y31, x0_y32, x1_y32, x2_y32, x3_y32, x4_y32, x5_y32, x6_y32, x7_y32, x8_y32, x9_y32, x10_y32, x11_y32, x12_y32, x13_y32, x14_y32, x15_y32, x16_y32, x17_y32, x18_y32, x19_y32, x20_y32, x21_y32, x22_y32, x23_y32, x24_y32, x25_y32, x26_y32, x27_y32, x28_y32, x29_y32, x30_y32, x31_y32, x32_y32, x33_y32, x34_y32, x35_y32, x36_y32, x37_y32, x38_y32, x39_y32, x40_y32, x41_y32, x42_y32, x43_y32, x44_y32, x45_y32, x46_y32, x47_y32, x48_y32, x0_y33, x1_y33, x2_y33, x3_y33, x4_y33, x5_y33, x6_y33, x7_y33, x8_y33, x9_y33, x10_y33, x11_y33, x12_y33, x13_y33, x14_y33, x15_y33, x16_y33, x17_y33, x18_y33, x19_y33, x20_y33, x21_y33, x22_y33, x23_y33, x24_y33, x25_y33, x26_y33, x27_y33, x28_y33, x29_y33, x30_y33, x31_y33, x32_y33, x33_y33, x34_y33, x35_y33, x36_y33, x37_y33, x38_y33, x39_y33, x40_y33, x41_y33, x42_y33, x43_y33, x44_y33, x45_y33, x46_y33, x47_y33, x48_y33, x0_y34, x1_y34, x2_y34, x3_y34, x4_y34, x5_y34, x6_y34, x7_y34, x8_y34, x9_y34, x10_y34, x11_y34, x12_y34, x13_y34, x14_y34, x15_y34, x16_y34, x17_y34, x18_y34, x19_y34, x20_y34, x21_y34, x22_y34, x23_y34, x24_y34, x25_y34, x26_y34, x27_y34, x28_y34, x29_y34, x30_y34, x31_y34, x32_y34, x33_y34, x34_y34, x35_y34, x36_y34, x37_y34, x38_y34, x39_y34, x40_y34, x41_y34, x42_y34, x43_y34, x44_y34, x45_y34, x46_y34, x47_y34, x48_y34, x0_y35, x1_y35, x2_y35, x3_y35, x4_y35, x5_y35, x6_y35, x7_y35, x8_y35, x9_y35, x10_y35, x11_y35, x12_y35, x13_y35, x14_y35, x15_y35, x16_y35, x17_y35, x18_y35, x19_y35, x20_y35, x21_y35, x22_y35, x23_y35, x24_y35, x25_y35, x26_y35, x27_y35, x28_y35, x29_y35, x30_y35, x31_y35, x32_y35, x33_y35, x34_y35, x35_y35, x36_y35, x37_y35, x38_y35, x39_y35, x40_y35, x41_y35, x42_y35, x43_y35, x44_y35, x45_y35, x46_y35, x47_y35, x48_y35, x0_y36, x1_y36, x2_y36, x3_y36, x4_y36, x5_y36, x6_y36, x7_y36, x8_y36, x9_y36, x10_y36, x11_y36, x12_y36, x13_y36, x14_y36, x15_y36, x16_y36, x17_y36, x18_y36, x19_y36, x20_y36, x21_y36, x22_y36, x23_y36, x24_y36, x25_y36, x26_y36, x27_y36, x28_y36, x29_y36, x30_y36, x31_y36, x32_y36, x33_y36, x34_y36, x35_y36, x36_y36, x37_y36, x38_y36, x39_y36, x40_y36, x41_y36, x42_y36, x43_y36, x44_y36, x45_y36, x46_y36, x47_y36, x48_y36, x0_y37, x1_y37, x2_y37, x3_y37, x4_y37, x5_y37, x6_y37, x7_y37, x8_y37, x9_y37, x10_y37, x11_y37, x12_y37, x13_y37, x14_y37, x15_y37, x16_y37, x17_y37, x18_y37, x19_y37, x20_y37, x21_y37, x22_y37, x23_y37, x24_y37, x25_y37, x26_y37, x27_y37, x28_y37, x29_y37, x30_y37, x31_y37, x32_y37, x33_y37, x34_y37, x35_y37, x36_y37, x37_y37, x38_y37, x39_y37, x40_y37, x41_y37, x42_y37, x43_y37, x44_y37, x45_y37, x46_y37, x47_y37, x48_y37, x0_y38, x1_y38, x2_y38, x3_y38, x4_y38, x5_y38, x6_y38, x7_y38, x8_y38, x9_y38, x10_y38, x11_y38, x12_y38, x13_y38, x14_y38, x15_y38, x16_y38, x17_y38, x18_y38, x19_y38, x20_y38, x21_y38, x22_y38, x23_y38, x24_y38, x25_y38, x26_y38, x27_y38, x28_y38, x29_y38, x30_y38, x31_y38, x32_y38, x33_y38, x34_y38, x35_y38, x36_y38, x37_y38, x38_y38, x39_y38, x40_y38, x41_y38, x42_y38, x43_y38, x44_y38, x45_y38, x46_y38, x47_y38, x48_y38, x0_y39, x1_y39, x2_y39, x3_y39, x4_y39, x5_y39, x6_y39, x7_y39, x8_y39, x9_y39, x10_y39, x11_y39, x12_y39, x13_y39, x14_y39, x15_y39, x16_y39, x17_y39, x18_y39, x19_y39, x20_y39, x21_y39, x22_y39, x23_y39, x24_y39, x25_y39, x26_y39, x27_y39, x28_y39, x29_y39, x30_y39, x31_y39, x32_y39, x33_y39, x34_y39, x35_y39, x36_y39, x37_y39, x38_y39, x39_y39, x40_y39, x41_y39, x42_y39, x43_y39, x44_y39, x45_y39, x46_y39, x47_y39, x48_y39, x0_y40, x1_y40, x2_y40, x3_y40, x4_y40, x5_y40, x6_y40, x7_y40, x8_y40, x9_y40, x10_y40, x11_y40, x12_y40, x13_y40, x14_y40, x15_y40, x16_y40, x17_y40, x18_y40, x19_y40, x20_y40, x21_y40, x22_y40, x23_y40, x24_y40, x25_y40, x26_y40, x27_y40, x28_y40, x29_y40, x30_y40, x31_y40, x32_y40, x33_y40, x34_y40, x35_y40, x36_y40, x37_y40, x38_y40, x39_y40, x40_y40, x41_y40, x42_y40, x43_y40, x44_y40, x45_y40, x46_y40, x47_y40, x48_y40, x0_y41, x1_y41, x2_y41, x3_y41, x4_y41, x5_y41, x6_y41, x7_y41, x8_y41, x9_y41, x10_y41, x11_y41, x12_y41, x13_y41, x14_y41, x15_y41, x16_y41, x17_y41, x18_y41, x19_y41, x20_y41, x21_y41, x22_y41, x23_y41, x24_y41, x25_y41, x26_y41, x27_y41, x28_y41, x29_y41, x30_y41, x31_y41, x32_y41, x33_y41, x34_y41, x35_y41, x36_y41, x37_y41, x38_y41, x39_y41, x40_y41, x41_y41, x42_y41, x43_y41, x44_y41, x45_y41, x46_y41, x47_y41, x48_y41, x0_y42, x1_y42, x2_y42, x3_y42, x4_y42, x5_y42, x6_y42, x7_y42, x8_y42, x9_y42, x10_y42, x11_y42, x12_y42, x13_y42, x14_y42, x15_y42, x16_y42, x17_y42, x18_y42, x19_y42, x20_y42, x21_y42, x22_y42, x23_y42, x24_y42, x25_y42, x26_y42, x27_y42, x28_y42, x29_y42, x30_y42, x31_y42, x32_y42, x33_y42, x34_y42, x35_y42, x36_y42, x37_y42, x38_y42, x39_y42, x40_y42, x41_y42, x42_y42, x43_y42, x44_y42, x45_y42, x46_y42, x47_y42, x48_y42, x0_y43, x1_y43, x2_y43, x3_y43, x4_y43, x5_y43, x6_y43, x7_y43, x8_y43, x9_y43, x10_y43, x11_y43, x12_y43, x13_y43, x14_y43, x15_y43, x16_y43, x17_y43, x18_y43, x19_y43, x20_y43, x21_y43, x22_y43, x23_y43, x24_y43, x25_y43, x26_y43, x27_y43, x28_y43, x29_y43, x30_y43, x31_y43, x32_y43, x33_y43, x34_y43, x35_y43, x36_y43, x37_y43, x38_y43, x39_y43, x40_y43, x41_y43, x42_y43, x43_y43, x44_y43, x45_y43, x46_y43, x47_y43, x48_y43, x0_y44, x1_y44, x2_y44, x3_y44, x4_y44, x5_y44, x6_y44, x7_y44, x8_y44, x9_y44, x10_y44, x11_y44, x12_y44, x13_y44, x14_y44, x15_y44, x16_y44, x17_y44, x18_y44, x19_y44, x20_y44, x21_y44, x22_y44, x23_y44, x24_y44, x25_y44, x26_y44, x27_y44, x28_y44, x29_y44, x30_y44, x31_y44, x32_y44, x33_y44, x34_y44, x35_y44, x36_y44, x37_y44, x38_y44, x39_y44, x40_y44, x41_y44, x42_y44, x43_y44, x44_y44, x45_y44, x46_y44, x47_y44, x48_y44, x0_y45, x1_y45, x2_y45, x3_y45, x4_y45, x5_y45, x6_y45, x7_y45, x8_y45, x9_y45, x10_y45, x11_y45, x12_y45, x13_y45, x14_y45, x15_y45, x16_y45, x17_y45, x18_y45, x19_y45, x20_y45, x21_y45, x22_y45, x23_y45, x24_y45, x25_y45, x26_y45, x27_y45, x28_y45, x29_y45, x30_y45, x31_y45, x32_y45, x33_y45, x34_y45, x35_y45, x36_y45, x37_y45, x38_y45, x39_y45, x40_y45, x41_y45, x42_y45, x43_y45, x44_y45, x45_y45, x46_y45, x47_y45, x48_y45, x0_y46, x1_y46, x2_y46, x3_y46, x4_y46, x5_y46, x6_y46, x7_y46, x8_y46, x9_y46, x10_y46, x11_y46, x12_y46, x13_y46, x14_y46, x15_y46, x16_y46, x17_y46, x18_y46, x19_y46, x20_y46, x21_y46, x22_y46, x23_y46, x24_y46, x25_y46, x26_y46, x27_y46, x28_y46, x29_y46, x30_y46, x31_y46, x32_y46, x33_y46, x34_y46, x35_y46, x36_y46, x37_y46, x38_y46, x39_y46, x40_y46, x41_y46, x42_y46, x43_y46, x44_y46, x45_y46, x46_y46, x47_y46, x48_y46, x0_y47, x1_y47, x2_y47, x3_y47, x4_y47, x5_y47, x6_y47, x7_y47, x8_y47, x9_y47, x10_y47, x11_y47, x12_y47, x13_y47, x14_y47, x15_y47, x16_y47, x17_y47, x18_y47, x19_y47, x20_y47, x21_y47, x22_y47, x23_y47, x24_y47, x25_y47, x26_y47, x27_y47, x28_y47, x29_y47, x30_y47, x31_y47, x32_y47, x33_y47, x34_y47, x35_y47, x36_y47, x37_y47, x38_y47, x39_y47, x40_y47, x41_y47, x42_y47, x43_y47, x44_y47, x45_y47, x46_y47, x47_y47, x48_y47, x0_y48, x1_y48, x2_y48, x3_y48, x4_y48, x5_y48, x6_y48, x7_y48, x8_y48, x9_y48, x10_y48, x11_y48, x12_y48, x13_y48, x14_y48, x15_y48, x16_y48, x17_y48, x18_y48, x19_y48, x20_y48, x21_y48, x22_y48, x23_y48, x24_y48, x25_y48, x26_y48, x27_y48, x28_y48, x29_y48, x30_y48, x31_y48, x32_y48, x33_y48, x34_y48, x35_y48, x36_y48, x37_y48, x38_y48, x39_y48, x40_y48, x41_y48, x42_y48, x43_y48, x44_y48, x45_y48, x46_y48, x47_y48, x48_y48, x0_y49, x1_y49, x2_y49, x3_y49, x4_y49, x5_y49, x6_y49, x7_y49, x8_y49, x9_y49, x10_y49, x11_y49, x12_y49, x13_y49, x14_y49, x15_y49, x16_y49, x17_y49, x18_y49, x19_y49, x20_y49, x21_y49, x22_y49, x23_y49, x24_y49, x25_y49, x26_y49, x27_y49, x28_y49, x29_y49, x30_y49, x31_y49, x32_y49, x33_y49, x34_y49, x35_y49, x36_y49, x37_y49, x38_y49, x39_y49, x40_y49, x41_y49, x42_y49, x43_y49, x44_y49, x45_y49, x46_y49, x47_y49, x48_y49;


(* keep, dont_touch *)
(* LOC = "X0/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011101101111)
) lut_0_0 (
    .O(x0_y0),
    .I0(in0),
    .I1(in2),
    .I2(in3),
    .I3(in0)
);

(* keep, dont_touch *)
(* LOC = "X1/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010000000000)
) lut_1_0 (
    .O(x1_y0),
    .I0(in4),
    .I1(1'b0),
    .I2(in0),
    .I3(in5)
);

(* keep, dont_touch *)
(* LOC = "X2/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001100010001)
) lut_2_0 (
    .O(x2_y0),
    .I0(1'b0),
    .I1(in1),
    .I2(in0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X3/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001001000111)
) lut_3_0 (
    .O(x3_y0),
    .I0(x1_y0),
    .I1(x1_y0),
    .I2(x1_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X4/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111100010111)
) lut_4_0 (
    .O(x4_y0),
    .I0(x2_y0),
    .I1(x1_y0),
    .I2(x2_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X5/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110000001010)
) lut_5_0 (
    .O(x5_y0),
    .I0(x2_y0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x2_y0)
);

(* keep, dont_touch *)
(* LOC = "X6/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001111111000)
) lut_6_0 (
    .O(x6_y0),
    .I0(x4_y4),
    .I1(x3_y0),
    .I2(x3_y0),
    .I3(x3_y1)
);

(* keep, dont_touch *)
(* LOC = "X7/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001111101101)
) lut_7_0 (
    .O(x7_y0),
    .I0(x5_y3),
    .I1(x4_y0),
    .I2(x4_y2),
    .I3(x5_y1)
);

(* keep, dont_touch *)
(* LOC = "X8/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111001101110)
) lut_8_0 (
    .O(x8_y0),
    .I0(x5_y0),
    .I1(x6_y0),
    .I2(x5_y0),
    .I3(x6_y0)
);

(* keep, dont_touch *)
(* LOC = "X9/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001010101110)
) lut_9_0 (
    .O(x9_y0),
    .I0(x6_y0),
    .I1(x6_y0),
    .I2(x5_y0),
    .I3(x6_y0)
);

(* keep, dont_touch *)
(* LOC = "X10/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101100111000)
) lut_10_0 (
    .O(x10_y0),
    .I0(1'b0),
    .I1(x8_y4),
    .I2(1'b0),
    .I3(x8_y5)
);

(* keep, dont_touch *)
(* LOC = "X11/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011000101100)
) lut_11_0 (
    .O(x11_y0),
    .I0(x9_y5),
    .I1(x8_y0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X12/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101101101011)
) lut_12_0 (
    .O(x12_y0),
    .I0(x10_y0),
    .I1(1'b0),
    .I2(x10_y5),
    .I3(x9_y0)
);

(* keep, dont_touch *)
(* LOC = "X13/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001011001111)
) lut_13_0 (
    .O(x13_y0),
    .I0(x11_y0),
    .I1(x10_y0),
    .I2(x11_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X14/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001111110011)
) lut_14_0 (
    .O(x14_y0),
    .I0(x11_y4),
    .I1(1'b0),
    .I2(x12_y5),
    .I3(x11_y5)
);

(* keep, dont_touch *)
(* LOC = "X15/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100101110100)
) lut_15_0 (
    .O(x15_y0),
    .I0(x12_y0),
    .I1(1'b0),
    .I2(x12_y0),
    .I3(x12_y0)
);

(* keep, dont_touch *)
(* LOC = "X16/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011010100101)
) lut_16_0 (
    .O(x16_y0),
    .I0(x13_y0),
    .I1(x13_y4),
    .I2(1'b0),
    .I3(x14_y0)
);

(* keep, dont_touch *)
(* LOC = "X17/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001101111010)
) lut_17_0 (
    .O(x17_y0),
    .I0(x15_y5),
    .I1(1'b0),
    .I2(x15_y0),
    .I3(x15_y0)
);

(* keep, dont_touch *)
(* LOC = "X18/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110000111111)
) lut_18_0 (
    .O(x18_y0),
    .I0(x16_y4),
    .I1(x15_y2),
    .I2(x15_y2),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X19/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100000111111)
) lut_19_0 (
    .O(x19_y0),
    .I0(x16_y1),
    .I1(1'b0),
    .I2(x16_y0),
    .I3(x16_y1)
);

(* keep, dont_touch *)
(* LOC = "X20/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000000000011)
) lut_20_0 (
    .O(x20_y0),
    .I0(x17_y3),
    .I1(x17_y0),
    .I2(x17_y1),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X21/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011010010100)
) lut_21_0 (
    .O(x21_y0),
    .I0(x18_y0),
    .I1(1'b0),
    .I2(x19_y0),
    .I3(x19_y4)
);

(* keep, dont_touch *)
(* LOC = "X22/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000111001111)
) lut_22_0 (
    .O(x22_y0),
    .I0(x19_y5),
    .I1(x20_y3),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X23/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110111011001)
) lut_23_0 (
    .O(x23_y0),
    .I0(x20_y2),
    .I1(x20_y0),
    .I2(x21_y5),
    .I3(x20_y4)
);

(* keep, dont_touch *)
(* LOC = "X24/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101000010111)
) lut_24_0 (
    .O(x24_y0),
    .I0(x22_y1),
    .I1(x22_y3),
    .I2(x22_y0),
    .I3(x22_y0)
);

(* keep, dont_touch *)
(* LOC = "X25/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100011111001)
) lut_25_0 (
    .O(x25_y0),
    .I0(x22_y0),
    .I1(x23_y0),
    .I2(x23_y0),
    .I3(x23_y3)
);

(* keep, dont_touch *)
(* LOC = "X26/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110010110111)
) lut_26_0 (
    .O(x26_y0),
    .I0(1'b0),
    .I1(x24_y3),
    .I2(x24_y3),
    .I3(x24_y5)
);

(* keep, dont_touch *)
(* LOC = "X27/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101010010111)
) lut_27_0 (
    .O(x27_y0),
    .I0(x24_y0),
    .I1(x24_y5),
    .I2(x25_y0),
    .I3(x24_y4)
);

(* keep, dont_touch *)
(* LOC = "X28/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010110110101)
) lut_28_0 (
    .O(x28_y0),
    .I0(x25_y2),
    .I1(1'b0),
    .I2(x25_y4),
    .I3(x26_y0)
);

(* keep, dont_touch *)
(* LOC = "X29/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011010100010)
) lut_29_0 (
    .O(x29_y0),
    .I0(x26_y0),
    .I1(x26_y5),
    .I2(x26_y0),
    .I3(x26_y3)
);

(* keep, dont_touch *)
(* LOC = "X30/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110100010111)
) lut_30_0 (
    .O(x30_y0),
    .I0(x27_y1),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x28_y0)
);

(* keep, dont_touch *)
(* LOC = "X31/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011011011010)
) lut_31_0 (
    .O(x31_y0),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x28_y3)
);

(* keep, dont_touch *)
(* LOC = "X32/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010101110100)
) lut_32_0 (
    .O(x32_y0),
    .I0(x30_y0),
    .I1(x29_y4),
    .I2(x30_y5),
    .I3(x29_y4)
);

(* keep, dont_touch *)
(* LOC = "X33/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101010111100)
) lut_33_0 (
    .O(x33_y0),
    .I0(1'b0),
    .I1(x30_y0),
    .I2(x30_y0),
    .I3(x30_y0)
);

(* keep, dont_touch *)
(* LOC = "X34/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000111010111)
) lut_34_0 (
    .O(x34_y0),
    .I0(x31_y3),
    .I1(x32_y0),
    .I2(x32_y0),
    .I3(x31_y3)
);

(* keep, dont_touch *)
(* LOC = "X35/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011110100010)
) lut_35_0 (
    .O(x35_y0),
    .I0(x32_y0),
    .I1(1'b0),
    .I2(x32_y2),
    .I3(x32_y0)
);

(* keep, dont_touch *)
(* LOC = "X36/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110110100110)
) lut_36_0 (
    .O(x36_y0),
    .I0(x33_y0),
    .I1(x34_y1),
    .I2(x33_y2),
    .I3(x34_y3)
);

(* keep, dont_touch *)
(* LOC = "X37/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000100001100)
) lut_37_0 (
    .O(x37_y0),
    .I0(1'b0),
    .I1(x34_y4),
    .I2(x35_y0),
    .I3(x35_y2)
);

(* keep, dont_touch *)
(* LOC = "X38/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011100110101)
) lut_38_0 (
    .O(x38_y0),
    .I0(x35_y3),
    .I1(x36_y3),
    .I2(x35_y2),
    .I3(x35_y0)
);

(* keep, dont_touch *)
(* LOC = "X39/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001110001001)
) lut_39_0 (
    .O(x39_y0),
    .I0(x36_y0),
    .I1(x37_y0),
    .I2(x36_y0),
    .I3(x37_y0)
);

(* keep, dont_touch *)
(* LOC = "X40/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001001110001)
) lut_40_0 (
    .O(x40_y0),
    .I0(1'b0),
    .I1(x37_y5),
    .I2(x37_y0),
    .I3(x37_y2)
);

(* keep, dont_touch *)
(* LOC = "X41/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100011010111)
) lut_41_0 (
    .O(x41_y0),
    .I0(x39_y0),
    .I1(x39_y0),
    .I2(x39_y0),
    .I3(x38_y0)
);

(* keep, dont_touch *)
(* LOC = "X42/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010100100001)
) lut_42_0 (
    .O(x42_y0),
    .I0(x39_y2),
    .I1(x39_y4),
    .I2(x39_y0),
    .I3(x40_y1)
);

(* keep, dont_touch *)
(* LOC = "X43/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000100111101)
) lut_43_0 (
    .O(x43_y0),
    .I0(x40_y1),
    .I1(x40_y2),
    .I2(1'b0),
    .I3(x40_y5)
);

(* keep, dont_touch *)
(* LOC = "X44/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100110101100)
) lut_44_0 (
    .O(x44_y0),
    .I0(x41_y0),
    .I1(1'b0),
    .I2(x41_y0),
    .I3(x41_y0)
);

(* keep, dont_touch *)
(* LOC = "X45/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011011100111)
) lut_45_0 (
    .O(x45_y0),
    .I0(x42_y0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x43_y0)
);

(* keep, dont_touch *)
(* LOC = "X46/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110000101110)
) lut_46_0 (
    .O(x46_y0),
    .I0(1'b0),
    .I1(x43_y5),
    .I2(1'b0),
    .I3(x43_y0)
);

(* keep, dont_touch *)
(* LOC = "X47/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010001100110)
) lut_47_0 (
    .O(x47_y0),
    .I0(x44_y3),
    .I1(x45_y0),
    .I2(x44_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X48/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010010000010)
) lut_48_0 (
    .O(x48_y0),
    .I0(1'b0),
    .I1(x46_y0),
    .I2(x46_y0),
    .I3(x46_y0)
);

(* keep, dont_touch *)
(* LOC = "X49/Y0" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100010100000)
) lut_49_0 (
    .O(x49_y0),
    .I0(x46_y2),
    .I1(x46_y0),
    .I2(x47_y0),
    .I3(x47_y0)
);

(* keep, dont_touch *)
(* LOC = "X0/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010110000000)
) lut_0_1 (
    .O(x0_y1),
    .I0(in0),
    .I1(in2),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X1/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101111101011)
) lut_1_1 (
    .O(x1_y1),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(in0)
);

(* keep, dont_touch *)
(* LOC = "X2/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001101000001)
) lut_2_1 (
    .O(x2_y1),
    .I0(in0),
    .I1(in4),
    .I2(in5),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X3/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111110101101)
) lut_3_1 (
    .O(x3_y1),
    .I0(x1_y2),
    .I1(x1_y1),
    .I2(1'b0),
    .I3(in0)
);

(* keep, dont_touch *)
(* LOC = "X4/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101100010110)
) lut_4_1 (
    .O(x4_y1),
    .I0(1'b0),
    .I1(x2_y0),
    .I2(x2_y5),
    .I3(x2_y0)
);

(* keep, dont_touch *)
(* LOC = "X5/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000010001111)
) lut_5_1 (
    .O(x5_y1),
    .I0(x2_y2),
    .I1(x2_y3),
    .I2(1'b0),
    .I3(x3_y0)
);

(* keep, dont_touch *)
(* LOC = "X6/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101100100001)
) lut_6_1 (
    .O(x6_y1),
    .I0(x3_y2),
    .I1(x3_y0),
    .I2(x4_y0),
    .I3(x4_y0)
);

(* keep, dont_touch *)
(* LOC = "X7/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111000001110)
) lut_7_1 (
    .O(x7_y1),
    .I0(x4_y2),
    .I1(x4_y2),
    .I2(x5_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X8/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001001011110)
) lut_8_1 (
    .O(x8_y1),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x6_y3),
    .I3(x6_y0)
);

(* keep, dont_touch *)
(* LOC = "X9/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101110101010)
) lut_9_1 (
    .O(x9_y1),
    .I0(x6_y6),
    .I1(x7_y5),
    .I2(x6_y3),
    .I3(x6_y0)
);

(* keep, dont_touch *)
(* LOC = "X10/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010000110001)
) lut_10_1 (
    .O(x10_y1),
    .I0(1'b0),
    .I1(x8_y0),
    .I2(1'b0),
    .I3(x7_y5)
);

(* keep, dont_touch *)
(* LOC = "X11/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110011101110)
) lut_11_1 (
    .O(x11_y1),
    .I0(x8_y3),
    .I1(x9_y1),
    .I2(x9_y0),
    .I3(x9_y0)
);

(* keep, dont_touch *)
(* LOC = "X12/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111110111110)
) lut_12_1 (
    .O(x12_y1),
    .I0(x9_y2),
    .I1(x9_y0),
    .I2(x10_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X13/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010110011000)
) lut_13_1 (
    .O(x13_y1),
    .I0(1'b0),
    .I1(x11_y4),
    .I2(x11_y4),
    .I3(x11_y4)
);

(* keep, dont_touch *)
(* LOC = "X14/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001010001100)
) lut_14_1 (
    .O(x14_y1),
    .I0(x12_y5),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X15/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110100111000)
) lut_15_1 (
    .O(x15_y1),
    .I0(1'b0),
    .I1(x13_y0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X16/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111101110011)
) lut_16_1 (
    .O(x16_y1),
    .I0(x13_y3),
    .I1(x14_y6),
    .I2(x13_y2),
    .I3(x13_y2)
);

(* keep, dont_touch *)
(* LOC = "X17/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100011001011)
) lut_17_1 (
    .O(x17_y1),
    .I0(x14_y5),
    .I1(x14_y5),
    .I2(1'b0),
    .I3(x15_y0)
);

(* keep, dont_touch *)
(* LOC = "X18/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110001010000)
) lut_18_1 (
    .O(x18_y1),
    .I0(x16_y3),
    .I1(x15_y0),
    .I2(x16_y0),
    .I3(x16_y1)
);

(* keep, dont_touch *)
(* LOC = "X19/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000011111011)
) lut_19_1 (
    .O(x19_y1),
    .I0(x16_y6),
    .I1(x16_y1),
    .I2(1'b0),
    .I3(x17_y0)
);

(* keep, dont_touch *)
(* LOC = "X20/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100100101001)
) lut_20_1 (
    .O(x20_y1),
    .I0(x18_y2),
    .I1(x18_y2),
    .I2(x17_y6),
    .I3(x18_y0)
);

(* keep, dont_touch *)
(* LOC = "X21/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110011101001)
) lut_21_1 (
    .O(x21_y1),
    .I0(x18_y5),
    .I1(1'b0),
    .I2(x19_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X22/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001101000101)
) lut_22_1 (
    .O(x22_y1),
    .I0(x20_y2),
    .I1(x19_y6),
    .I2(1'b0),
    .I3(x20_y2)
);

(* keep, dont_touch *)
(* LOC = "X23/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011001101001)
) lut_23_1 (
    .O(x23_y1),
    .I0(x21_y3),
    .I1(x21_y2),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X24/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111001100101)
) lut_24_1 (
    .O(x24_y1),
    .I0(x22_y6),
    .I1(x21_y4),
    .I2(1'b0),
    .I3(x22_y4)
);

(* keep, dont_touch *)
(* LOC = "X25/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100101100100)
) lut_25_1 (
    .O(x25_y1),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x22_y6),
    .I3(x23_y0)
);

(* keep, dont_touch *)
(* LOC = "X26/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001010110110)
) lut_26_1 (
    .O(x26_y1),
    .I0(x23_y0),
    .I1(1'b0),
    .I2(x24_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X27/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010011001001)
) lut_27_1 (
    .O(x27_y1),
    .I0(x25_y0),
    .I1(1'b0),
    .I2(x24_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X28/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111000100101)
) lut_28_1 (
    .O(x28_y1),
    .I0(x26_y0),
    .I1(1'b0),
    .I2(x25_y1),
    .I3(x25_y0)
);

(* keep, dont_touch *)
(* LOC = "X29/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010101011111)
) lut_29_1 (
    .O(x29_y1),
    .I0(x26_y0),
    .I1(x26_y3),
    .I2(x26_y6),
    .I3(x26_y1)
);

(* keep, dont_touch *)
(* LOC = "X30/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000111100101)
) lut_30_1 (
    .O(x30_y1),
    .I0(x27_y0),
    .I1(x27_y0),
    .I2(1'b0),
    .I3(x27_y0)
);

(* keep, dont_touch *)
(* LOC = "X31/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100010011100)
) lut_31_1 (
    .O(x31_y1),
    .I0(1'b0),
    .I1(x29_y5),
    .I2(x29_y0),
    .I3(x28_y0)
);

(* keep, dont_touch *)
(* LOC = "X32/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011100110110)
) lut_32_1 (
    .O(x32_y1),
    .I0(x30_y0),
    .I1(x29_y0),
    .I2(x29_y5),
    .I3(x30_y2)
);

(* keep, dont_touch *)
(* LOC = "X33/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101000110110)
) lut_33_1 (
    .O(x33_y1),
    .I0(x31_y4),
    .I1(1'b0),
    .I2(x30_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X34/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110111000111)
) lut_34_1 (
    .O(x34_y1),
    .I0(x31_y1),
    .I1(x32_y0),
    .I2(x31_y0),
    .I3(x31_y0)
);

(* keep, dont_touch *)
(* LOC = "X35/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011101011001)
) lut_35_1 (
    .O(x35_y1),
    .I0(x32_y0),
    .I1(x32_y3),
    .I2(x32_y3),
    .I3(x32_y4)
);

(* keep, dont_touch *)
(* LOC = "X36/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000110101011)
) lut_36_1 (
    .O(x36_y1),
    .I0(1'b0),
    .I1(x34_y0),
    .I2(x33_y2),
    .I3(x33_y0)
);

(* keep, dont_touch *)
(* LOC = "X37/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001011011011)
) lut_37_1 (
    .O(x37_y1),
    .I0(x34_y1),
    .I1(x35_y0),
    .I2(1'b0),
    .I3(x35_y0)
);

(* keep, dont_touch *)
(* LOC = "X38/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000011101011)
) lut_38_1 (
    .O(x38_y1),
    .I0(x35_y2),
    .I1(x36_y1),
    .I2(x35_y1),
    .I3(x36_y6)
);

(* keep, dont_touch *)
(* LOC = "X39/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111011101101)
) lut_39_1 (
    .O(x39_y1),
    .I0(x37_y0),
    .I1(x36_y0),
    .I2(x37_y6),
    .I3(x37_y1)
);

(* keep, dont_touch *)
(* LOC = "X40/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100110101000)
) lut_40_1 (
    .O(x40_y1),
    .I0(x38_y0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x37_y0)
);

(* keep, dont_touch *)
(* LOC = "X41/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011110101010)
) lut_41_1 (
    .O(x41_y1),
    .I0(1'b0),
    .I1(x38_y1),
    .I2(x38_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X42/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100111010100)
) lut_42_1 (
    .O(x42_y1),
    .I0(x39_y2),
    .I1(x40_y2),
    .I2(x39_y3),
    .I3(x39_y6)
);

(* keep, dont_touch *)
(* LOC = "X43/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101010101111)
) lut_43_1 (
    .O(x43_y1),
    .I0(x40_y5),
    .I1(x40_y4),
    .I2(x40_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X44/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010010111111)
) lut_44_1 (
    .O(x44_y1),
    .I0(x42_y2),
    .I1(x41_y0),
    .I2(x41_y1),
    .I3(x41_y0)
);

(* keep, dont_touch *)
(* LOC = "X45/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011110110001)
) lut_45_1 (
    .O(x45_y1),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X46/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101111111101)
) lut_46_1 (
    .O(x46_y1),
    .I0(x44_y1),
    .I1(1'b0),
    .I2(x44_y3),
    .I3(x43_y0)
);

(* keep, dont_touch *)
(* LOC = "X47/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001100110111)
) lut_47_1 (
    .O(x47_y1),
    .I0(1'b0),
    .I1(x45_y0),
    .I2(x44_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X48/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101100011110)
) lut_48_1 (
    .O(x48_y1),
    .I0(x46_y1),
    .I1(x46_y4),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X49/Y1" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000101010100)
) lut_49_1 (
    .O(x49_y1),
    .I0(x47_y0),
    .I1(x46_y0),
    .I2(x47_y4),
    .I3(x47_y0)
);

(* keep, dont_touch *)
(* LOC = "X0/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010101110100)
) lut_0_2 (
    .O(x0_y2),
    .I0(1'b0),
    .I1(in2),
    .I2(in5),
    .I3(in5)
);

(* keep, dont_touch *)
(* LOC = "X1/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110010001111)
) lut_1_2 (
    .O(x1_y2),
    .I0(in5),
    .I1(in0),
    .I2(1'b0),
    .I3(in7)
);

(* keep, dont_touch *)
(* LOC = "X2/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001110100010)
) lut_2_2 (
    .O(x2_y2),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X3/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110110101001)
) lut_3_2 (
    .O(x3_y2),
    .I0(1'b0),
    .I1(in5),
    .I2(x1_y6),
    .I3(x1_y4)
);

(* keep, dont_touch *)
(* LOC = "X4/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101110110011)
) lut_4_2 (
    .O(x4_y2),
    .I0(x1_y2),
    .I1(x2_y3),
    .I2(x1_y4),
    .I3(x1_y7)
);

(* keep, dont_touch *)
(* LOC = "X5/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010001011001)
) lut_5_2 (
    .O(x5_y2),
    .I0(x2_y0),
    .I1(x2_y3),
    .I2(x2_y2),
    .I3(x3_y4)
);

(* keep, dont_touch *)
(* LOC = "X6/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100011101100)
) lut_6_2 (
    .O(x6_y2),
    .I0(x3_y0),
    .I1(x3_y0),
    .I2(x4_y4),
    .I3(x3_y0)
);

(* keep, dont_touch *)
(* LOC = "X7/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001010111101)
) lut_7_2 (
    .O(x7_y2),
    .I0(1'b0),
    .I1(x4_y0),
    .I2(x5_y0),
    .I3(x5_y0)
);

(* keep, dont_touch *)
(* LOC = "X8/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100100111110)
) lut_8_2 (
    .O(x8_y2),
    .I0(x5_y0),
    .I1(x6_y0),
    .I2(x6_y0),
    .I3(x5_y3)
);

(* keep, dont_touch *)
(* LOC = "X9/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001011101011)
) lut_9_2 (
    .O(x9_y2),
    .I0(x7_y0),
    .I1(1'b0),
    .I2(x6_y0),
    .I3(x5_y3)
);

(* keep, dont_touch *)
(* LOC = "X10/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110000001111)
) lut_10_2 (
    .O(x10_y2),
    .I0(x8_y0),
    .I1(1'b0),
    .I2(x7_y4),
    .I3(x7_y2)
);

(* keep, dont_touch *)
(* LOC = "X11/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010010110011)
) lut_11_2 (
    .O(x11_y2),
    .I0(x9_y0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X12/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000100110101)
) lut_12_2 (
    .O(x12_y2),
    .I0(x9_y3),
    .I1(x9_y4),
    .I2(x9_y1),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X13/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101001011111)
) lut_13_2 (
    .O(x13_y2),
    .I0(x10_y2),
    .I1(x10_y1),
    .I2(x10_y1),
    .I3(x10_y3)
);

(* keep, dont_touch *)
(* LOC = "X14/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011011101000)
) lut_14_2 (
    .O(x14_y2),
    .I0(x12_y1),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x11_y0)
);

(* keep, dont_touch *)
(* LOC = "X15/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001111111111)
) lut_15_2 (
    .O(x15_y2),
    .I0(x12_y3),
    .I1(x13_y5),
    .I2(x13_y2),
    .I3(x13_y3)
);

(* keep, dont_touch *)
(* LOC = "X16/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110000101111)
) lut_16_2 (
    .O(x16_y2),
    .I0(x13_y0),
    .I1(x14_y2),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X17/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000000000010)
) lut_17_2 (
    .O(x17_y2),
    .I0(x15_y0),
    .I1(x14_y5),
    .I2(1'b0),
    .I3(x14_y2)
);

(* keep, dont_touch *)
(* LOC = "X18/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111011110010)
) lut_18_2 (
    .O(x18_y2),
    .I0(1'b0),
    .I1(x16_y0),
    .I2(x16_y0),
    .I3(x16_y5)
);

(* keep, dont_touch *)
(* LOC = "X19/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000001110111)
) lut_19_2 (
    .O(x19_y2),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x17_y7),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X20/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100000010001)
) lut_20_2 (
    .O(x20_y2),
    .I0(x17_y2),
    .I1(1'b0),
    .I2(x18_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X21/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101110010111)
) lut_21_2 (
    .O(x21_y2),
    .I0(x18_y0),
    .I1(1'b0),
    .I2(x18_y0),
    .I3(x19_y0)
);

(* keep, dont_touch *)
(* LOC = "X22/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010001110010)
) lut_22_2 (
    .O(x22_y2),
    .I0(x20_y5),
    .I1(x20_y6),
    .I2(1'b0),
    .I3(x19_y0)
);

(* keep, dont_touch *)
(* LOC = "X23/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011111001100)
) lut_23_2 (
    .O(x23_y2),
    .I0(1'b0),
    .I1(x21_y0),
    .I2(x20_y7),
    .I3(x20_y7)
);

(* keep, dont_touch *)
(* LOC = "X24/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001000000100)
) lut_24_2 (
    .O(x24_y2),
    .I0(x21_y1),
    .I1(1'b0),
    .I2(x21_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X25/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011101000110)
) lut_25_2 (
    .O(x25_y2),
    .I0(x22_y0),
    .I1(x22_y1),
    .I2(x23_y0),
    .I3(x23_y3)
);

(* keep, dont_touch *)
(* LOC = "X26/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010110010110)
) lut_26_2 (
    .O(x26_y2),
    .I0(x24_y0),
    .I1(x24_y6),
    .I2(x24_y1),
    .I3(x24_y6)
);

(* keep, dont_touch *)
(* LOC = "X27/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010000100110)
) lut_27_2 (
    .O(x27_y2),
    .I0(x24_y0),
    .I1(x25_y0),
    .I2(x25_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X28/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001000110011)
) lut_28_2 (
    .O(x28_y2),
    .I0(x26_y0),
    .I1(x26_y3),
    .I2(1'b0),
    .I3(x26_y0)
);

(* keep, dont_touch *)
(* LOC = "X29/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011111000100)
) lut_29_2 (
    .O(x29_y2),
    .I0(x26_y5),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x26_y7)
);

(* keep, dont_touch *)
(* LOC = "X30/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101000011010)
) lut_30_2 (
    .O(x30_y2),
    .I0(x27_y0),
    .I1(x27_y4),
    .I2(x28_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X31/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101000100010)
) lut_31_2 (
    .O(x31_y2),
    .I0(x29_y0),
    .I1(x29_y1),
    .I2(x29_y7),
    .I3(x28_y6)
);

(* keep, dont_touch *)
(* LOC = "X32/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110001010110)
) lut_32_2 (
    .O(x32_y2),
    .I0(x29_y1),
    .I1(x30_y0),
    .I2(x30_y0),
    .I3(x30_y1)
);

(* keep, dont_touch *)
(* LOC = "X33/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001010000101)
) lut_33_2 (
    .O(x33_y2),
    .I0(x31_y0),
    .I1(x31_y7),
    .I2(x31_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X34/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110010110110)
) lut_34_2 (
    .O(x34_y2),
    .I0(1'b0),
    .I1(x31_y3),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X35/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101110100100)
) lut_35_2 (
    .O(x35_y2),
    .I0(1'b0),
    .I1(x32_y7),
    .I2(1'b0),
    .I3(x33_y1)
);

(* keep, dont_touch *)
(* LOC = "X36/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110101010111)
) lut_36_2 (
    .O(x36_y2),
    .I0(x33_y5),
    .I1(x34_y5),
    .I2(x33_y0),
    .I3(x34_y0)
);

(* keep, dont_touch *)
(* LOC = "X37/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101101111101)
) lut_37_2 (
    .O(x37_y2),
    .I0(x34_y0),
    .I1(1'b0),
    .I2(x34_y5),
    .I3(x34_y5)
);

(* keep, dont_touch *)
(* LOC = "X38/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100010111000)
) lut_38_2 (
    .O(x38_y2),
    .I0(x35_y0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x35_y2)
);

(* keep, dont_touch *)
(* LOC = "X39/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111111010100)
) lut_39_2 (
    .O(x39_y2),
    .I0(x36_y0),
    .I1(x37_y3),
    .I2(x36_y6),
    .I3(x36_y7)
);

(* keep, dont_touch *)
(* LOC = "X40/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011010010010)
) lut_40_2 (
    .O(x40_y2),
    .I0(x38_y2),
    .I1(x38_y2),
    .I2(1'b0),
    .I3(x38_y5)
);

(* keep, dont_touch *)
(* LOC = "X41/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011110011001)
) lut_41_2 (
    .O(x41_y2),
    .I0(x38_y2),
    .I1(x38_y0),
    .I2(x39_y0),
    .I3(x38_y2)
);

(* keep, dont_touch *)
(* LOC = "X42/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100101001101)
) lut_42_2 (
    .O(x42_y2),
    .I0(x40_y0),
    .I1(x39_y0),
    .I2(1'b0),
    .I3(x39_y6)
);

(* keep, dont_touch *)
(* LOC = "X43/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010110101110)
) lut_43_2 (
    .O(x43_y2),
    .I0(x40_y4),
    .I1(x41_y0),
    .I2(x41_y0),
    .I3(x40_y1)
);

(* keep, dont_touch *)
(* LOC = "X44/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100011111100)
) lut_44_2 (
    .O(x44_y2),
    .I0(1'b0),
    .I1(x41_y4),
    .I2(x41_y0),
    .I3(x41_y0)
);

(* keep, dont_touch *)
(* LOC = "X45/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001001000001)
) lut_45_2 (
    .O(x45_y2),
    .I0(x43_y0),
    .I1(x42_y0),
    .I2(x43_y1),
    .I3(x42_y4)
);

(* keep, dont_touch *)
(* LOC = "X46/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111100101101)
) lut_46_2 (
    .O(x46_y2),
    .I0(x43_y3),
    .I1(x43_y6),
    .I2(x44_y4),
    .I3(x44_y7)
);

(* keep, dont_touch *)
(* LOC = "X47/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000000110000)
) lut_47_2 (
    .O(x47_y2),
    .I0(x44_y2),
    .I1(x45_y2),
    .I2(x44_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X48/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111101000001)
) lut_48_2 (
    .O(x48_y2),
    .I0(1'b0),
    .I1(x45_y2),
    .I2(x46_y6),
    .I3(x46_y7)
);

(* keep, dont_touch *)
(* LOC = "X49/Y2" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001111000101)
) lut_49_2 (
    .O(x49_y2),
    .I0(x47_y5),
    .I1(x46_y0),
    .I2(x46_y0),
    .I3(x47_y0)
);

(* keep, dont_touch *)
(* LOC = "X0/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101011000010)
) lut_0_3 (
    .O(x0_y3),
    .I0(in0),
    .I1(in2),
    .I2(in0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X1/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101100100000)
) lut_1_3 (
    .O(x1_y3),
    .I0(in0),
    .I1(1'b0),
    .I2(in3),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X2/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101110000111)
) lut_2_3 (
    .O(x2_y3),
    .I0(1'b0),
    .I1(in7),
    .I2(1'b0),
    .I3(in4)
);

(* keep, dont_touch *)
(* LOC = "X3/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111000111100)
) lut_3_3 (
    .O(x3_y3),
    .I0(in2),
    .I1(1'b0),
    .I2(1'b0),
    .I3(in1)
);

(* keep, dont_touch *)
(* LOC = "X4/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100111001011)
) lut_4_3 (
    .O(x4_y3),
    .I0(x1_y0),
    .I1(x2_y5),
    .I2(1'b0),
    .I3(x2_y1)
);

(* keep, dont_touch *)
(* LOC = "X5/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011100111110)
) lut_5_3 (
    .O(x5_y3),
    .I0(x3_y0),
    .I1(x3_y1),
    .I2(x3_y0),
    .I3(x3_y5)
);

(* keep, dont_touch *)
(* LOC = "X6/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110110011010)
) lut_6_3 (
    .O(x6_y3),
    .I0(1'b0),
    .I1(x4_y6),
    .I2(x3_y3),
    .I3(x3_y1)
);

(* keep, dont_touch *)
(* LOC = "X7/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011010011000)
) lut_7_3 (
    .O(x7_y3),
    .I0(x4_y0),
    .I1(1'b0),
    .I2(x4_y7),
    .I3(x5_y1)
);

(* keep, dont_touch *)
(* LOC = "X8/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000111110110)
) lut_8_3 (
    .O(x8_y3),
    .I0(1'b0),
    .I1(x6_y4),
    .I2(x6_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X9/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010010100001)
) lut_9_3 (
    .O(x9_y3),
    .I0(1'b0),
    .I1(x7_y5),
    .I2(x6_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X10/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001101011111)
) lut_10_3 (
    .O(x10_y3),
    .I0(x7_y8),
    .I1(1'b0),
    .I2(x7_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X11/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000100010001)
) lut_11_3 (
    .O(x11_y3),
    .I0(x9_y0),
    .I1(x8_y0),
    .I2(x8_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X12/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000101011010)
) lut_12_3 (
    .O(x12_y3),
    .I0(1'b0),
    .I1(x10_y8),
    .I2(x10_y0),
    .I3(x9_y0)
);

(* keep, dont_touch *)
(* LOC = "X13/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000111101001)
) lut_13_3 (
    .O(x13_y3),
    .I0(x10_y1),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x10_y3)
);

(* keep, dont_touch *)
(* LOC = "X14/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001000011010)
) lut_14_3 (
    .O(x14_y3),
    .I0(x11_y3),
    .I1(1'b0),
    .I2(x11_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X15/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101001101110)
) lut_15_3 (
    .O(x15_y3),
    .I0(x12_y1),
    .I1(x13_y4),
    .I2(x12_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X16/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111001000011)
) lut_16_3 (
    .O(x16_y3),
    .I0(x14_y0),
    .I1(1'b0),
    .I2(x13_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X17/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011011100110)
) lut_17_3 (
    .O(x17_y3),
    .I0(1'b0),
    .I1(x15_y0),
    .I2(x14_y2),
    .I3(x15_y1)
);

(* keep, dont_touch *)
(* LOC = "X18/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010100001111)
) lut_18_3 (
    .O(x18_y3),
    .I0(1'b0),
    .I1(x15_y3),
    .I2(x15_y0),
    .I3(x15_y3)
);

(* keep, dont_touch *)
(* LOC = "X19/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111110101010)
) lut_19_3 (
    .O(x19_y3),
    .I0(x16_y7),
    .I1(1'b0),
    .I2(x17_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X20/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010101110001)
) lut_20_3 (
    .O(x20_y3),
    .I0(x18_y1),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x18_y1)
);

(* keep, dont_touch *)
(* LOC = "X21/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111011111001)
) lut_21_3 (
    .O(x21_y3),
    .I0(x18_y2),
    .I1(1'b0),
    .I2(x18_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X22/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101110100001)
) lut_22_3 (
    .O(x22_y3),
    .I0(1'b0),
    .I1(x20_y1),
    .I2(x20_y0),
    .I3(x19_y3)
);

(* keep, dont_touch *)
(* LOC = "X23/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110100111010)
) lut_23_3 (
    .O(x23_y3),
    .I0(x20_y3),
    .I1(x20_y2),
    .I2(x21_y6),
    .I3(x21_y8)
);

(* keep, dont_touch *)
(* LOC = "X24/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111111011101)
) lut_24_3 (
    .O(x24_y3),
    .I0(x21_y6),
    .I1(x21_y6),
    .I2(x21_y4),
    .I3(x22_y4)
);

(* keep, dont_touch *)
(* LOC = "X25/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111110001101)
) lut_25_3 (
    .O(x25_y3),
    .I0(1'b0),
    .I1(x23_y2),
    .I2(x23_y5),
    .I3(x23_y3)
);

(* keep, dont_touch *)
(* LOC = "X26/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111111010110)
) lut_26_3 (
    .O(x26_y3),
    .I0(x23_y6),
    .I1(x24_y6),
    .I2(x23_y2),
    .I3(x24_y6)
);

(* keep, dont_touch *)
(* LOC = "X27/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111101101001)
) lut_27_3 (
    .O(x27_y3),
    .I0(x24_y4),
    .I1(x24_y2),
    .I2(x24_y0),
    .I3(x25_y1)
);

(* keep, dont_touch *)
(* LOC = "X28/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001010010011)
) lut_28_3 (
    .O(x28_y3),
    .I0(1'b0),
    .I1(x25_y3),
    .I2(1'b0),
    .I3(x26_y5)
);

(* keep, dont_touch *)
(* LOC = "X29/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011111110010)
) lut_29_3 (
    .O(x29_y3),
    .I0(1'b0),
    .I1(x27_y0),
    .I2(x26_y6),
    .I3(x26_y8)
);

(* keep, dont_touch *)
(* LOC = "X30/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001100010110)
) lut_30_3 (
    .O(x30_y3),
    .I0(x27_y7),
    .I1(x28_y0),
    .I2(1'b0),
    .I3(x28_y3)
);

(* keep, dont_touch *)
(* LOC = "X31/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100000100100)
) lut_31_3 (
    .O(x31_y3),
    .I0(1'b0),
    .I1(x29_y8),
    .I2(x28_y7),
    .I3(x28_y8)
);

(* keep, dont_touch *)
(* LOC = "X32/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010111010010)
) lut_32_3 (
    .O(x32_y3),
    .I0(x29_y5),
    .I1(x30_y4),
    .I2(x30_y5),
    .I3(x29_y0)
);

(* keep, dont_touch *)
(* LOC = "X33/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010010010001)
) lut_33_3 (
    .O(x33_y3),
    .I0(x30_y0),
    .I1(x31_y7),
    .I2(x30_y5),
    .I3(x30_y1)
);

(* keep, dont_touch *)
(* LOC = "X34/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011011000010)
) lut_34_3 (
    .O(x34_y3),
    .I0(x31_y6),
    .I1(x31_y0),
    .I2(1'b0),
    .I3(x32_y4)
);

(* keep, dont_touch *)
(* LOC = "X35/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101101001101)
) lut_35_3 (
    .O(x35_y3),
    .I0(x32_y6),
    .I1(x33_y0),
    .I2(x32_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X36/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001111101011)
) lut_36_3 (
    .O(x36_y3),
    .I0(x34_y8),
    .I1(x34_y6),
    .I2(x34_y0),
    .I3(x33_y3)
);

(* keep, dont_touch *)
(* LOC = "X37/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010111111100)
) lut_37_3 (
    .O(x37_y3),
    .I0(x34_y0),
    .I1(1'b0),
    .I2(x34_y2),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X38/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100101101000)
) lut_38_3 (
    .O(x38_y3),
    .I0(x36_y2),
    .I1(x35_y1),
    .I2(x36_y0),
    .I3(x36_y6)
);

(* keep, dont_touch *)
(* LOC = "X39/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000110001010)
) lut_39_3 (
    .O(x39_y3),
    .I0(x37_y0),
    .I1(1'b0),
    .I2(x36_y1),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X40/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001000011000)
) lut_40_3 (
    .O(x40_y3),
    .I0(1'b0),
    .I1(x38_y0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X41/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100011100000)
) lut_41_3 (
    .O(x41_y3),
    .I0(x38_y2),
    .I1(x38_y0),
    .I2(x38_y6),
    .I3(x38_y4)
);

(* keep, dont_touch *)
(* LOC = "X42/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111111000010)
) lut_42_3 (
    .O(x42_y3),
    .I0(x40_y5),
    .I1(x40_y6),
    .I2(x39_y6),
    .I3(x40_y0)
);

(* keep, dont_touch *)
(* LOC = "X43/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101110001011)
) lut_43_3 (
    .O(x43_y3),
    .I0(x40_y4),
    .I1(1'b0),
    .I2(x40_y1),
    .I3(x41_y4)
);

(* keep, dont_touch *)
(* LOC = "X44/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101100011111)
) lut_44_3 (
    .O(x44_y3),
    .I0(x41_y8),
    .I1(x42_y0),
    .I2(x42_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X45/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111110110100)
) lut_45_3 (
    .O(x45_y3),
    .I0(x43_y0),
    .I1(x42_y0),
    .I2(x42_y4),
    .I3(x42_y2)
);

(* keep, dont_touch *)
(* LOC = "X46/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010100101010)
) lut_46_3 (
    .O(x46_y3),
    .I0(x44_y6),
    .I1(x44_y8),
    .I2(x43_y3),
    .I3(x43_y4)
);

(* keep, dont_touch *)
(* LOC = "X47/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000011100111)
) lut_47_3 (
    .O(x47_y3),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x44_y2),
    .I3(x45_y7)
);

(* keep, dont_touch *)
(* LOC = "X48/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111000101000)
) lut_48_3 (
    .O(x48_y3),
    .I0(x46_y0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x46_y4)
);

(* keep, dont_touch *)
(* LOC = "X49/Y3" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010000001011)
) lut_49_3 (
    .O(x49_y3),
    .I0(x47_y0),
    .I1(x46_y8),
    .I2(x46_y4),
    .I3(x46_y5)
);

(* keep, dont_touch *)
(* LOC = "X0/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011110101010)
) lut_0_4 (
    .O(x0_y4),
    .I0(1'b0),
    .I1(in4),
    .I2(in3),
    .I3(in7)
);

(* keep, dont_touch *)
(* LOC = "X1/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010010010101)
) lut_1_4 (
    .O(x1_y4),
    .I0(in1),
    .I1(in1),
    .I2(in8),
    .I3(in3)
);

(* keep, dont_touch *)
(* LOC = "X2/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100001011000)
) lut_2_4 (
    .O(x2_y4),
    .I0(in3),
    .I1(in8),
    .I2(in6),
    .I3(in4)
);

(* keep, dont_touch *)
(* LOC = "X3/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111100010011)
) lut_3_4 (
    .O(x3_y4),
    .I0(x1_y0),
    .I1(in2),
    .I2(in7),
    .I3(in0)
);

(* keep, dont_touch *)
(* LOC = "X4/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001101101111)
) lut_4_4 (
    .O(x4_y4),
    .I0(x2_y1),
    .I1(x2_y0),
    .I2(x1_y7),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X5/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110100000100)
) lut_5_4 (
    .O(x5_y4),
    .I0(x2_y8),
    .I1(x2_y0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X6/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010000010000)
) lut_6_4 (
    .O(x6_y4),
    .I0(1'b0),
    .I1(x3_y2),
    .I2(x3_y2),
    .I3(x3_y3)
);

(* keep, dont_touch *)
(* LOC = "X7/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111010110010)
) lut_7_4 (
    .O(x7_y4),
    .I0(1'b0),
    .I1(x5_y3),
    .I2(x5_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X8/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101000001100)
) lut_8_4 (
    .O(x8_y4),
    .I0(x6_y1),
    .I1(x5_y2),
    .I2(x5_y4),
    .I3(x5_y0)
);

(* keep, dont_touch *)
(* LOC = "X9/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000110100000)
) lut_9_4 (
    .O(x9_y4),
    .I0(x7_y1),
    .I1(x7_y8),
    .I2(x5_y4),
    .I3(x5_y0)
);

(* keep, dont_touch *)
(* LOC = "X10/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011100101010)
) lut_10_4 (
    .O(x10_y4),
    .I0(x7_y9),
    .I1(x7_y7),
    .I2(x7_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X11/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000011110000)
) lut_11_4 (
    .O(x11_y4),
    .I0(1'b0),
    .I1(x9_y1),
    .I2(x9_y1),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X12/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110101111010)
) lut_12_4 (
    .O(x12_y4),
    .I0(x9_y5),
    .I1(x10_y2),
    .I2(x10_y8),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X13/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010100010011)
) lut_13_4 (
    .O(x13_y4),
    .I0(x11_y0),
    .I1(x11_y3),
    .I2(x10_y1),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X14/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100001110111)
) lut_14_4 (
    .O(x14_y4),
    .I0(x11_y9),
    .I1(x11_y1),
    .I2(1'b0),
    .I3(x11_y9)
);

(* keep, dont_touch *)
(* LOC = "X15/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100010100110)
) lut_15_4 (
    .O(x15_y4),
    .I0(1'b0),
    .I1(x13_y0),
    .I2(x12_y2),
    .I3(x12_y1)
);

(* keep, dont_touch *)
(* LOC = "X16/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010011001111)
) lut_16_4 (
    .O(x16_y4),
    .I0(x13_y9),
    .I1(x13_y0),
    .I2(x14_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X17/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010000111001)
) lut_17_4 (
    .O(x17_y4),
    .I0(x14_y2),
    .I1(x14_y9),
    .I2(x15_y8),
    .I3(x14_y5)
);

(* keep, dont_touch *)
(* LOC = "X18/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101111000111)
) lut_18_4 (
    .O(x18_y4),
    .I0(x16_y7),
    .I1(x15_y1),
    .I2(x15_y2),
    .I3(x15_y0)
);

(* keep, dont_touch *)
(* LOC = "X19/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110110100111)
) lut_19_4 (
    .O(x19_y4),
    .I0(x16_y0),
    .I1(x17_y7),
    .I2(x17_y0),
    .I3(x17_y5)
);

(* keep, dont_touch *)
(* LOC = "X20/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101101100010)
) lut_20_4 (
    .O(x20_y4),
    .I0(x18_y6),
    .I1(x17_y8),
    .I2(1'b0),
    .I3(x17_y5)
);

(* keep, dont_touch *)
(* LOC = "X21/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111011101000)
) lut_21_4 (
    .O(x21_y4),
    .I0(x18_y8),
    .I1(1'b0),
    .I2(x19_y1),
    .I3(x18_y0)
);

(* keep, dont_touch *)
(* LOC = "X22/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101100110111)
) lut_22_4 (
    .O(x22_y4),
    .I0(x20_y5),
    .I1(x19_y9),
    .I2(x20_y5),
    .I3(x19_y6)
);

(* keep, dont_touch *)
(* LOC = "X23/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100100110111)
) lut_23_4 (
    .O(x23_y4),
    .I0(x21_y5),
    .I1(1'b0),
    .I2(x21_y6),
    .I3(x21_y4)
);

(* keep, dont_touch *)
(* LOC = "X24/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011110101110)
) lut_24_4 (
    .O(x24_y4),
    .I0(1'b0),
    .I1(x21_y5),
    .I2(x22_y0),
    .I3(x22_y0)
);

(* keep, dont_touch *)
(* LOC = "X25/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000001011101)
) lut_25_4 (
    .O(x25_y4),
    .I0(x22_y7),
    .I1(x23_y0),
    .I2(x23_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X26/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001011010001)
) lut_26_4 (
    .O(x26_y4),
    .I0(x23_y1),
    .I1(x24_y4),
    .I2(x24_y2),
    .I3(x24_y7)
);

(* keep, dont_touch *)
(* LOC = "X27/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100011010101)
) lut_27_4 (
    .O(x27_y4),
    .I0(x24_y4),
    .I1(x24_y0),
    .I2(1'b0),
    .I3(x24_y1)
);

(* keep, dont_touch *)
(* LOC = "X28/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100000001110)
) lut_28_4 (
    .O(x28_y4),
    .I0(x26_y8),
    .I1(x25_y0),
    .I2(x26_y0),
    .I3(x26_y6)
);

(* keep, dont_touch *)
(* LOC = "X29/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010111110111)
) lut_29_4 (
    .O(x29_y4),
    .I0(x27_y7),
    .I1(x26_y2),
    .I2(x26_y0),
    .I3(x27_y7)
);

(* keep, dont_touch *)
(* LOC = "X30/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001010001011)
) lut_30_4 (
    .O(x30_y4),
    .I0(x28_y0),
    .I1(x27_y6),
    .I2(1'b0),
    .I3(x27_y3)
);

(* keep, dont_touch *)
(* LOC = "X31/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111011100010)
) lut_31_4 (
    .O(x31_y4),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x28_y6)
);

(* keep, dont_touch *)
(* LOC = "X32/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110000000011)
) lut_32_4 (
    .O(x32_y4),
    .I0(x30_y9),
    .I1(x30_y4),
    .I2(x30_y0),
    .I3(x29_y6)
);

(* keep, dont_touch *)
(* LOC = "X33/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110000001100)
) lut_33_4 (
    .O(x33_y4),
    .I0(x31_y6),
    .I1(x30_y0),
    .I2(x31_y9),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X34/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110000110100)
) lut_34_4 (
    .O(x34_y4),
    .I0(x32_y1),
    .I1(x32_y4),
    .I2(x32_y3),
    .I3(x32_y6)
);

(* keep, dont_touch *)
(* LOC = "X35/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100101101100)
) lut_35_4 (
    .O(x35_y4),
    .I0(x33_y5),
    .I1(1'b0),
    .I2(x32_y0),
    .I3(x32_y4)
);

(* keep, dont_touch *)
(* LOC = "X36/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011100101101)
) lut_36_4 (
    .O(x36_y4),
    .I0(1'b0),
    .I1(x33_y0),
    .I2(1'b0),
    .I3(x34_y9)
);

(* keep, dont_touch *)
(* LOC = "X37/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000101001110)
) lut_37_4 (
    .O(x37_y4),
    .I0(x34_y0),
    .I1(1'b0),
    .I2(x34_y9),
    .I3(x35_y0)
);

(* keep, dont_touch *)
(* LOC = "X38/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101101101101)
) lut_38_4 (
    .O(x38_y4),
    .I0(x36_y4),
    .I1(x35_y1),
    .I2(x36_y9),
    .I3(x36_y4)
);

(* keep, dont_touch *)
(* LOC = "X39/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001101111001)
) lut_39_4 (
    .O(x39_y4),
    .I0(x36_y0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x37_y0)
);

(* keep, dont_touch *)
(* LOC = "X40/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111001001011)
) lut_40_4 (
    .O(x40_y4),
    .I0(x38_y4),
    .I1(x37_y3),
    .I2(x38_y4),
    .I3(x37_y4)
);

(* keep, dont_touch *)
(* LOC = "X41/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011000110101)
) lut_41_4 (
    .O(x41_y4),
    .I0(1'b0),
    .I1(x38_y3),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X42/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010111001111)
) lut_42_4 (
    .O(x42_y4),
    .I0(x40_y0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X43/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111000010001)
) lut_43_4 (
    .O(x43_y4),
    .I0(x41_y3),
    .I1(x41_y5),
    .I2(1'b0),
    .I3(x40_y1)
);

(* keep, dont_touch *)
(* LOC = "X44/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100001100101)
) lut_44_4 (
    .O(x44_y4),
    .I0(x42_y0),
    .I1(1'b0),
    .I2(x41_y7),
    .I3(x41_y0)
);

(* keep, dont_touch *)
(* LOC = "X45/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010001100000)
) lut_45_4 (
    .O(x45_y4),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x43_y7)
);

(* keep, dont_touch *)
(* LOC = "X46/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011000000110)
) lut_46_4 (
    .O(x46_y4),
    .I0(x43_y8),
    .I1(1'b0),
    .I2(x44_y0),
    .I3(x43_y6)
);

(* keep, dont_touch *)
(* LOC = "X47/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011000101101)
) lut_47_4 (
    .O(x47_y4),
    .I0(x45_y6),
    .I1(x44_y4),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X48/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101111001110)
) lut_48_4 (
    .O(x48_y4),
    .I0(x46_y8),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x46_y0)
);

(* keep, dont_touch *)
(* LOC = "X49/Y4" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110011001111)
) lut_49_4 (
    .O(x49_y4),
    .I0(x47_y1),
    .I1(x46_y9),
    .I2(x46_y7),
    .I3(x46_y0)
);

(* keep, dont_touch *)
(* LOC = "X0/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101111100011)
) lut_0_5 (
    .O(x0_y5),
    .I0(in7),
    .I1(in3),
    .I2(in9),
    .I3(in3)
);

(* keep, dont_touch *)
(* LOC = "X1/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011100010110)
) lut_1_5 (
    .O(x1_y5),
    .I0(in5),
    .I1(1'b0),
    .I2(in2),
    .I3(in4)
);

(* keep, dont_touch *)
(* LOC = "X2/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101010011110)
) lut_2_5 (
    .O(x2_y5),
    .I0(in9),
    .I1(in2),
    .I2(in2),
    .I3(in0)
);

(* keep, dont_touch *)
(* LOC = "X3/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011010110001)
) lut_3_5 (
    .O(x3_y5),
    .I0(x1_y2),
    .I1(in0),
    .I2(1'b0),
    .I3(in0)
);

(* keep, dont_touch *)
(* LOC = "X4/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000111100110)
) lut_4_5 (
    .O(x4_y5),
    .I0(1'b0),
    .I1(x1_y5),
    .I2(x2_y6),
    .I3(x1_y10)
);

(* keep, dont_touch *)
(* LOC = "X5/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111101001110)
) lut_5_5 (
    .O(x5_y5),
    .I0(x2_y9),
    .I1(x2_y6),
    .I2(x2_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X6/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010100100110)
) lut_6_5 (
    .O(x6_y5),
    .I0(x4_y7),
    .I1(x4_y5),
    .I2(x3_y6),
    .I3(x3_y0)
);

(* keep, dont_touch *)
(* LOC = "X7/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100001101100)
) lut_7_5 (
    .O(x7_y5),
    .I0(1'b0),
    .I1(x4_y2),
    .I2(1'b0),
    .I3(x5_y3)
);

(* keep, dont_touch *)
(* LOC = "X8/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000101110101)
) lut_8_5 (
    .O(x8_y5),
    .I0(x5_y0),
    .I1(x5_y8),
    .I2(1'b0),
    .I3(x5_y7)
);

(* keep, dont_touch *)
(* LOC = "X9/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010111110111)
) lut_9_5 (
    .O(x9_y5),
    .I0(1'b0),
    .I1(x6_y4),
    .I2(1'b0),
    .I3(x5_y7)
);

(* keep, dont_touch *)
(* LOC = "X10/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011001110101)
) lut_10_5 (
    .O(x10_y5),
    .I0(x7_y1),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x8_y5)
);

(* keep, dont_touch *)
(* LOC = "X11/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001000111111)
) lut_11_5 (
    .O(x11_y5),
    .I0(x8_y7),
    .I1(x9_y6),
    .I2(x8_y2),
    .I3(x8_y2)
);

(* keep, dont_touch *)
(* LOC = "X12/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101101011011)
) lut_12_5 (
    .O(x12_y5),
    .I0(x9_y9),
    .I1(1'b0),
    .I2(x9_y2),
    .I3(x10_y4)
);

(* keep, dont_touch *)
(* LOC = "X13/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110010000101)
) lut_13_5 (
    .O(x13_y5),
    .I0(x10_y9),
    .I1(x11_y2),
    .I2(x11_y1),
    .I3(x11_y10)
);

(* keep, dont_touch *)
(* LOC = "X14/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000010100001)
) lut_14_5 (
    .O(x14_y5),
    .I0(x11_y3),
    .I1(x11_y9),
    .I2(x11_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X15/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111110000011)
) lut_15_5 (
    .O(x15_y5),
    .I0(1'b0),
    .I1(x13_y3),
    .I2(x12_y9),
    .I3(x13_y6)
);

(* keep, dont_touch *)
(* LOC = "X16/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000001110011)
) lut_16_5 (
    .O(x16_y5),
    .I0(x13_y5),
    .I1(x14_y3),
    .I2(x14_y1),
    .I3(x14_y7)
);

(* keep, dont_touch *)
(* LOC = "X17/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100111110100)
) lut_17_5 (
    .O(x17_y5),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x14_y7),
    .I3(x15_y5)
);

(* keep, dont_touch *)
(* LOC = "X18/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111010011110)
) lut_18_5 (
    .O(x18_y5),
    .I0(x16_y4),
    .I1(x16_y9),
    .I2(x16_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X19/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101010001000)
) lut_19_5 (
    .O(x19_y5),
    .I0(x16_y8),
    .I1(1'b0),
    .I2(x17_y5),
    .I3(x17_y9)
);

(* keep, dont_touch *)
(* LOC = "X20/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011111111001)
) lut_20_5 (
    .O(x20_y5),
    .I0(x18_y4),
    .I1(x17_y2),
    .I2(x17_y0),
    .I3(x17_y10)
);

(* keep, dont_touch *)
(* LOC = "X21/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010110110100)
) lut_21_5 (
    .O(x21_y5),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x19_y2),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X22/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110000011111)
) lut_22_5 (
    .O(x22_y5),
    .I0(x20_y8),
    .I1(x20_y3),
    .I2(x20_y7),
    .I3(x19_y4)
);

(* keep, dont_touch *)
(* LOC = "X23/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011011011010)
) lut_23_5 (
    .O(x23_y5),
    .I0(x20_y10),
    .I1(x20_y3),
    .I2(x21_y10),
    .I3(x21_y0)
);

(* keep, dont_touch *)
(* LOC = "X24/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010100000000)
) lut_24_5 (
    .O(x24_y5),
    .I0(x21_y9),
    .I1(1'b0),
    .I2(x22_y2),
    .I3(x22_y5)
);

(* keep, dont_touch *)
(* LOC = "X25/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000001000100)
) lut_25_5 (
    .O(x25_y5),
    .I0(x23_y7),
    .I1(1'b0),
    .I2(x23_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X26/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011110101100)
) lut_26_5 (
    .O(x26_y5),
    .I0(x24_y1),
    .I1(x24_y2),
    .I2(x23_y0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X27/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110000010100)
) lut_27_5 (
    .O(x27_y5),
    .I0(x24_y4),
    .I1(x24_y4),
    .I2(x24_y10),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X28/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111010100001)
) lut_28_5 (
    .O(x28_y5),
    .I0(x26_y7),
    .I1(1'b0),
    .I2(x25_y7),
    .I3(x25_y9)
);

(* keep, dont_touch *)
(* LOC = "X29/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100100110010)
) lut_29_5 (
    .O(x29_y5),
    .I0(1'b0),
    .I1(x27_y10),
    .I2(x27_y1),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X30/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111000010011)
) lut_30_5 (
    .O(x30_y5),
    .I0(x28_y1),
    .I1(x28_y2),
    .I2(x28_y5),
    .I3(x28_y7)
);

(* keep, dont_touch *)
(* LOC = "X31/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010111000010)
) lut_31_5 (
    .O(x31_y5),
    .I0(x28_y9),
    .I1(x28_y8),
    .I2(x28_y4),
    .I3(x28_y1)
);

(* keep, dont_touch *)
(* LOC = "X32/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101110001111)
) lut_32_5 (
    .O(x32_y5),
    .I0(x29_y5),
    .I1(x29_y4),
    .I2(x29_y7),
    .I3(x29_y2)
);

(* keep, dont_touch *)
(* LOC = "X33/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101010001001)
) lut_33_5 (
    .O(x33_y5),
    .I0(x31_y4),
    .I1(x30_y10),
    .I2(x31_y9),
    .I3(x30_y4)
);

(* keep, dont_touch *)
(* LOC = "X34/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100101010010)
) lut_34_5 (
    .O(x34_y5),
    .I0(x31_y6),
    .I1(x32_y0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X35/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010101111010)
) lut_35_5 (
    .O(x35_y5),
    .I0(x32_y2),
    .I1(x33_y1),
    .I2(x32_y7),
    .I3(x33_y10)
);

(* keep, dont_touch *)
(* LOC = "X36/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101110101011)
) lut_36_5 (
    .O(x36_y5),
    .I0(x33_y4),
    .I1(x34_y8),
    .I2(1'b0),
    .I3(x33_y2)
);

(* keep, dont_touch *)
(* LOC = "X37/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010101101000)
) lut_37_5 (
    .O(x37_y5),
    .I0(x35_y2),
    .I1(x34_y5),
    .I2(x35_y7),
    .I3(x34_y1)
);

(* keep, dont_touch *)
(* LOC = "X38/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101001100010)
) lut_38_5 (
    .O(x38_y5),
    .I0(x35_y9),
    .I1(x36_y10),
    .I2(x36_y5),
    .I3(x35_y7)
);

(* keep, dont_touch *)
(* LOC = "X39/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001110110100)
) lut_39_5 (
    .O(x39_y5),
    .I0(1'b0),
    .I1(x36_y5),
    .I2(1'b0),
    .I3(x37_y1)
);

(* keep, dont_touch *)
(* LOC = "X40/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001010001010)
) lut_40_5 (
    .O(x40_y5),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x37_y9),
    .I3(x38_y4)
);

(* keep, dont_touch *)
(* LOC = "X41/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000101010000)
) lut_41_5 (
    .O(x41_y5),
    .I0(x38_y9),
    .I1(1'b0),
    .I2(x39_y1),
    .I3(x38_y4)
);

(* keep, dont_touch *)
(* LOC = "X42/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001111111111)
) lut_42_5 (
    .O(x42_y5),
    .I0(x40_y9),
    .I1(x40_y10),
    .I2(1'b0),
    .I3(x40_y1)
);

(* keep, dont_touch *)
(* LOC = "X43/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011111100100)
) lut_43_5 (
    .O(x43_y5),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x40_y6),
    .I3(x40_y9)
);

(* keep, dont_touch *)
(* LOC = "X44/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110011110011)
) lut_44_5 (
    .O(x44_y5),
    .I0(x41_y3),
    .I1(1'b0),
    .I2(x41_y3),
    .I3(x41_y6)
);

(* keep, dont_touch *)
(* LOC = "X45/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110000101101)
) lut_45_5 (
    .O(x45_y5),
    .I0(1'b0),
    .I1(x42_y3),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X46/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000011110111)
) lut_46_5 (
    .O(x46_y5),
    .I0(1'b0),
    .I1(x44_y3),
    .I2(1'b0),
    .I3(x43_y4)
);

(* keep, dont_touch *)
(* LOC = "X47/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101101011011)
) lut_47_5 (
    .O(x47_y5),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x45_y3),
    .I3(x45_y8)
);

(* keep, dont_touch *)
(* LOC = "X48/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010000101100)
) lut_48_5 (
    .O(x48_y5),
    .I0(x46_y4),
    .I1(x45_y6),
    .I2(x45_y6),
    .I3(x45_y0)
);

(* keep, dont_touch *)
(* LOC = "X49/Y5" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000001011010)
) lut_49_5 (
    .O(x49_y5),
    .I0(x46_y8),
    .I1(1'b0),
    .I2(x46_y8),
    .I3(x46_y1)
);

(* keep, dont_touch *)
(* LOC = "X0/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000001110000)
) lut_0_6 (
    .O(x0_y6),
    .I0(in4),
    .I1(1'b0),
    .I2(in5),
    .I3(in9)
);

(* keep, dont_touch *)
(* LOC = "X1/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010010010101)
) lut_1_6 (
    .O(x1_y6),
    .I0(in1),
    .I1(in9),
    .I2(in1),
    .I3(in8)
);

(* keep, dont_touch *)
(* LOC = "X2/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111010101001)
) lut_2_6 (
    .O(x2_y6),
    .I0(in8),
    .I1(in9),
    .I2(1'b0),
    .I3(in6)
);

(* keep, dont_touch *)
(* LOC = "X3/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110010000100)
) lut_3_6 (
    .O(x3_y6),
    .I0(x1_y1),
    .I1(in4),
    .I2(1'b0),
    .I3(in1)
);

(* keep, dont_touch *)
(* LOC = "X4/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011100000000)
) lut_4_6 (
    .O(x4_y6),
    .I0(x1_y2),
    .I1(x1_y7),
    .I2(1'b0),
    .I3(x1_y3)
);

(* keep, dont_touch *)
(* LOC = "X5/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001110010100)
) lut_5_6 (
    .O(x5_y6),
    .I0(x3_y3),
    .I1(x2_y4),
    .I2(x3_y9),
    .I3(x3_y8)
);

(* keep, dont_touch *)
(* LOC = "X6/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000000110101)
) lut_6_6 (
    .O(x6_y6),
    .I0(x4_y7),
    .I1(x3_y6),
    .I2(x3_y10),
    .I3(x3_y3)
);

(* keep, dont_touch *)
(* LOC = "X7/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110010001101)
) lut_7_6 (
    .O(x7_y6),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x4_y7)
);

(* keep, dont_touch *)
(* LOC = "X8/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011000101100)
) lut_8_6 (
    .O(x8_y6),
    .I0(1'b0),
    .I1(x5_y11),
    .I2(x6_y7),
    .I3(x5_y9)
);

(* keep, dont_touch *)
(* LOC = "X9/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101111100110)
) lut_9_6 (
    .O(x9_y6),
    .I0(x7_y3),
    .I1(1'b0),
    .I2(x6_y7),
    .I3(x5_y9)
);

(* keep, dont_touch *)
(* LOC = "X10/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011001010110)
) lut_10_6 (
    .O(x10_y6),
    .I0(x7_y2),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x7_y10)
);

(* keep, dont_touch *)
(* LOC = "X11/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001001101110)
) lut_11_6 (
    .O(x11_y6),
    .I0(x8_y7),
    .I1(x9_y6),
    .I2(x9_y9),
    .I3(x8_y10)
);

(* keep, dont_touch *)
(* LOC = "X12/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101110010000)
) lut_12_6 (
    .O(x12_y6),
    .I0(x9_y4),
    .I1(x9_y4),
    .I2(x10_y8),
    .I3(x9_y6)
);

(* keep, dont_touch *)
(* LOC = "X13/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110011001111)
) lut_13_6 (
    .O(x13_y6),
    .I0(x11_y1),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X14/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001100100110)
) lut_14_6 (
    .O(x14_y6),
    .I0(x11_y4),
    .I1(1'b0),
    .I2(x11_y5),
    .I3(x12_y10)
);

(* keep, dont_touch *)
(* LOC = "X15/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010010011111)
) lut_15_6 (
    .O(x15_y6),
    .I0(x12_y1),
    .I1(1'b0),
    .I2(x12_y1),
    .I3(x13_y3)
);

(* keep, dont_touch *)
(* LOC = "X16/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101111110001)
) lut_16_6 (
    .O(x16_y6),
    .I0(1'b0),
    .I1(x13_y6),
    .I2(x13_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X17/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111101001010)
) lut_17_6 (
    .O(x17_y6),
    .I0(x15_y5),
    .I1(x14_y5),
    .I2(x14_y1),
    .I3(x15_y4)
);

(* keep, dont_touch *)
(* LOC = "X18/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001101010000)
) lut_18_6 (
    .O(x18_y6),
    .I0(x15_y3),
    .I1(1'b0),
    .I2(x16_y4),
    .I3(x15_y1)
);

(* keep, dont_touch *)
(* LOC = "X19/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111100011011)
) lut_19_6 (
    .O(x19_y6),
    .I0(x16_y5),
    .I1(x17_y6),
    .I2(x17_y10),
    .I3(x17_y2)
);

(* keep, dont_touch *)
(* LOC = "X20/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001101101111)
) lut_20_6 (
    .O(x20_y6),
    .I0(x17_y3),
    .I1(x18_y6),
    .I2(x17_y10),
    .I3(x18_y1)
);

(* keep, dont_touch *)
(* LOC = "X21/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001100010010)
) lut_21_6 (
    .O(x21_y6),
    .I0(x19_y4),
    .I1(x18_y4),
    .I2(1'b0),
    .I3(x18_y9)
);

(* keep, dont_touch *)
(* LOC = "X22/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100100110000)
) lut_22_6 (
    .O(x22_y6),
    .I0(x19_y1),
    .I1(x19_y4),
    .I2(x20_y5),
    .I3(x19_y1)
);

(* keep, dont_touch *)
(* LOC = "X23/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010001110000)
) lut_23_6 (
    .O(x23_y6),
    .I0(1'b0),
    .I1(x20_y8),
    .I2(1'b0),
    .I3(x21_y11)
);

(* keep, dont_touch *)
(* LOC = "X24/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011101001110)
) lut_24_6 (
    .O(x24_y6),
    .I0(x21_y7),
    .I1(1'b0),
    .I2(x22_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X25/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100010001000)
) lut_25_6 (
    .O(x25_y6),
    .I0(x22_y9),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x23_y11)
);

(* keep, dont_touch *)
(* LOC = "X26/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110000100001)
) lut_26_6 (
    .O(x26_y6),
    .I0(x23_y8),
    .I1(x24_y11),
    .I2(x24_y5),
    .I3(x24_y6)
);

(* keep, dont_touch *)
(* LOC = "X27/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011101000111)
) lut_27_6 (
    .O(x27_y6),
    .I0(x25_y11),
    .I1(1'b0),
    .I2(x24_y2),
    .I3(x25_y5)
);

(* keep, dont_touch *)
(* LOC = "X28/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001111100111)
) lut_28_6 (
    .O(x28_y6),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x26_y6),
    .I3(x25_y7)
);

(* keep, dont_touch *)
(* LOC = "X29/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000001010111)
) lut_29_6 (
    .O(x29_y6),
    .I0(x26_y3),
    .I1(x27_y1),
    .I2(x27_y1),
    .I3(x27_y3)
);

(* keep, dont_touch *)
(* LOC = "X30/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001100011010)
) lut_30_6 (
    .O(x30_y6),
    .I0(x28_y4),
    .I1(x28_y5),
    .I2(1'b0),
    .I3(x27_y11)
);

(* keep, dont_touch *)
(* LOC = "X31/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100110110010)
) lut_31_6 (
    .O(x31_y6),
    .I0(x29_y11),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x29_y6)
);

(* keep, dont_touch *)
(* LOC = "X32/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001010101010)
) lut_32_6 (
    .O(x32_y6),
    .I0(x30_y7),
    .I1(x30_y3),
    .I2(x30_y5),
    .I3(x29_y6)
);

(* keep, dont_touch *)
(* LOC = "X33/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101101000100)
) lut_33_6 (
    .O(x33_y6),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x30_y4),
    .I3(x30_y10)
);

(* keep, dont_touch *)
(* LOC = "X34/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000010110100)
) lut_34_6 (
    .O(x34_y6),
    .I0(x31_y2),
    .I1(1'b0),
    .I2(x32_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X35/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001010001001)
) lut_35_6 (
    .O(x35_y6),
    .I0(1'b0),
    .I1(x32_y7),
    .I2(1'b0),
    .I3(x32_y7)
);

(* keep, dont_touch *)
(* LOC = "X36/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110101001101)
) lut_36_6 (
    .O(x36_y6),
    .I0(1'b0),
    .I1(x34_y10),
    .I2(x33_y4),
    .I3(x34_y4)
);

(* keep, dont_touch *)
(* LOC = "X37/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111001101000)
) lut_37_6 (
    .O(x37_y6),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x35_y2),
    .I3(x35_y8)
);

(* keep, dont_touch *)
(* LOC = "X38/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001101110011)
) lut_38_6 (
    .O(x38_y6),
    .I0(x36_y11),
    .I1(1'b0),
    .I2(x35_y5),
    .I3(x36_y1)
);

(* keep, dont_touch *)
(* LOC = "X39/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110011011010)
) lut_39_6 (
    .O(x39_y6),
    .I0(x37_y4),
    .I1(x37_y5),
    .I2(x37_y2),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X40/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001101001011)
) lut_40_6 (
    .O(x40_y6),
    .I0(x37_y6),
    .I1(x38_y10),
    .I2(x37_y6),
    .I3(x37_y4)
);

(* keep, dont_touch *)
(* LOC = "X41/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011110000010)
) lut_41_6 (
    .O(x41_y6),
    .I0(x39_y7),
    .I1(x38_y6),
    .I2(x38_y6),
    .I3(x39_y6)
);

(* keep, dont_touch *)
(* LOC = "X42/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010001001111)
) lut_42_6 (
    .O(x42_y6),
    .I0(x39_y4),
    .I1(x39_y6),
    .I2(x40_y6),
    .I3(x40_y11)
);

(* keep, dont_touch *)
(* LOC = "X43/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111000010011)
) lut_43_6 (
    .O(x43_y6),
    .I0(x40_y5),
    .I1(x41_y10),
    .I2(1'b0),
    .I3(x40_y2)
);

(* keep, dont_touch *)
(* LOC = "X44/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000001001100)
) lut_44_6 (
    .O(x44_y6),
    .I0(x42_y1),
    .I1(x42_y4),
    .I2(x41_y7),
    .I3(x41_y8)
);

(* keep, dont_touch *)
(* LOC = "X45/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000000111110)
) lut_45_6 (
    .O(x45_y6),
    .I0(x42_y8),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x43_y5)
);

(* keep, dont_touch *)
(* LOC = "X46/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110111001011)
) lut_46_6 (
    .O(x46_y6),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x44_y8),
    .I3(x44_y4)
);

(* keep, dont_touch *)
(* LOC = "X47/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011001011001)
) lut_47_6 (
    .O(x47_y6),
    .I0(1'b0),
    .I1(x45_y11),
    .I2(x45_y10),
    .I3(x44_y7)
);

(* keep, dont_touch *)
(* LOC = "X48/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110110000111)
) lut_48_6 (
    .O(x48_y6),
    .I0(x46_y7),
    .I1(x45_y2),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X49/Y6" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100001101111)
) lut_49_6 (
    .O(x49_y6),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x46_y5),
    .I3(x47_y2)
);

(* keep, dont_touch *)
(* LOC = "X0/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000011100111)
) lut_0_7 (
    .O(x0_y7),
    .I0(in1),
    .I1(in3),
    .I2(in3),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X1/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111011010000)
) lut_1_7 (
    .O(x1_y7),
    .I0(1'b0),
    .I1(in7),
    .I2(in5),
    .I3(in8)
);

(* keep, dont_touch *)
(* LOC = "X2/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001001100111)
) lut_2_7 (
    .O(x2_y7),
    .I0(in6),
    .I1(in2),
    .I2(in2),
    .I3(in6)
);

(* keep, dont_touch *)
(* LOC = "X3/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101001100000)
) lut_3_7 (
    .O(x3_y7),
    .I0(in5),
    .I1(1'b0),
    .I2(in5),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X4/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101110100000)
) lut_4_7 (
    .O(x4_y7),
    .I0(x2_y6),
    .I1(x1_y12),
    .I2(1'b0),
    .I3(x1_y8)
);

(* keep, dont_touch *)
(* LOC = "X5/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010001101100)
) lut_5_7 (
    .O(x5_y7),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x2_y3)
);

(* keep, dont_touch *)
(* LOC = "X6/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101100010100)
) lut_6_7 (
    .O(x6_y7),
    .I0(x3_y7),
    .I1(1'b0),
    .I2(x3_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X7/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100010100010)
) lut_7_7 (
    .O(x7_y7),
    .I0(x4_y9),
    .I1(x4_y7),
    .I2(x5_y12),
    .I3(x4_y4)
);

(* keep, dont_touch *)
(* LOC = "X8/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100011101100)
) lut_8_7 (
    .O(x8_y7),
    .I0(x6_y12),
    .I1(1'b0),
    .I2(x6_y10),
    .I3(x6_y3)
);

(* keep, dont_touch *)
(* LOC = "X9/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101110101101)
) lut_9_7 (
    .O(x9_y7),
    .I0(1'b0),
    .I1(x7_y4),
    .I2(x6_y10),
    .I3(x6_y3)
);

(* keep, dont_touch *)
(* LOC = "X10/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110100110001)
) lut_10_7 (
    .O(x10_y7),
    .I0(x8_y4),
    .I1(x8_y8),
    .I2(1'b0),
    .I3(x8_y10)
);

(* keep, dont_touch *)
(* LOC = "X11/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111010100000)
) lut_11_7 (
    .O(x11_y7),
    .I0(x9_y2),
    .I1(x9_y6),
    .I2(x8_y5),
    .I3(x9_y12)
);

(* keep, dont_touch *)
(* LOC = "X12/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110010000011)
) lut_12_7 (
    .O(x12_y7),
    .I0(1'b0),
    .I1(x9_y12),
    .I2(1'b0),
    .I3(x10_y11)
);

(* keep, dont_touch *)
(* LOC = "X13/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101110001001)
) lut_13_7 (
    .O(x13_y7),
    .I0(x11_y8),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x11_y12)
);

(* keep, dont_touch *)
(* LOC = "X14/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001001010000)
) lut_14_7 (
    .O(x14_y7),
    .I0(x11_y7),
    .I1(x11_y11),
    .I2(1'b0),
    .I3(x11_y4)
);

(* keep, dont_touch *)
(* LOC = "X15/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010011101001)
) lut_15_7 (
    .O(x15_y7),
    .I0(x13_y3),
    .I1(1'b0),
    .I2(x12_y11),
    .I3(x13_y12)
);

(* keep, dont_touch *)
(* LOC = "X16/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100010101100)
) lut_16_7 (
    .O(x16_y7),
    .I0(1'b0),
    .I1(x14_y7),
    .I2(x14_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X17/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110111100000)
) lut_17_7 (
    .O(x17_y7),
    .I0(x15_y10),
    .I1(x15_y11),
    .I2(x14_y11),
    .I3(x15_y10)
);

(* keep, dont_touch *)
(* LOC = "X18/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000110110110)
) lut_18_7 (
    .O(x18_y7),
    .I0(x15_y6),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x16_y4)
);

(* keep, dont_touch *)
(* LOC = "X19/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101011111111)
) lut_19_7 (
    .O(x19_y7),
    .I0(x17_y7),
    .I1(x16_y8),
    .I2(x16_y4),
    .I3(x17_y10)
);

(* keep, dont_touch *)
(* LOC = "X20/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110000110100)
) lut_20_7 (
    .O(x20_y7),
    .I0(1'b0),
    .I1(x17_y5),
    .I2(x17_y7),
    .I3(x18_y8)
);

(* keep, dont_touch *)
(* LOC = "X21/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101010011101)
) lut_21_7 (
    .O(x21_y7),
    .I0(x19_y2),
    .I1(x19_y6),
    .I2(x18_y4),
    .I3(x18_y6)
);

(* keep, dont_touch *)
(* LOC = "X22/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101110100110)
) lut_22_7 (
    .O(x22_y7),
    .I0(x20_y8),
    .I1(x19_y11),
    .I2(x20_y5),
    .I3(x20_y7)
);

(* keep, dont_touch *)
(* LOC = "X23/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110100110010)
) lut_23_7 (
    .O(x23_y7),
    .I0(x21_y6),
    .I1(x21_y9),
    .I2(x20_y12),
    .I3(x21_y6)
);

(* keep, dont_touch *)
(* LOC = "X24/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000110110100)
) lut_24_7 (
    .O(x24_y7),
    .I0(1'b0),
    .I1(x22_y8),
    .I2(x22_y2),
    .I3(x22_y3)
);

(* keep, dont_touch *)
(* LOC = "X25/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000011001101)
) lut_25_7 (
    .O(x25_y7),
    .I0(x23_y6),
    .I1(x23_y7),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X26/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000000000100)
) lut_26_7 (
    .O(x26_y7),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x24_y10),
    .I3(x24_y7)
);

(* keep, dont_touch *)
(* LOC = "X27/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001001110000)
) lut_27_7 (
    .O(x27_y7),
    .I0(1'b0),
    .I1(x24_y2),
    .I2(x24_y3),
    .I3(x25_y3)
);

(* keep, dont_touch *)
(* LOC = "X28/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101010000001)
) lut_28_7 (
    .O(x28_y7),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x26_y3),
    .I3(x26_y11)
);

(* keep, dont_touch *)
(* LOC = "X29/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111111111111)
) lut_29_7 (
    .O(x29_y7),
    .I0(x26_y12),
    .I1(x26_y8),
    .I2(x27_y8),
    .I3(x27_y5)
);

(* keep, dont_touch *)
(* LOC = "X30/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001111111100)
) lut_30_7 (
    .O(x30_y7),
    .I0(x28_y6),
    .I1(x27_y3),
    .I2(x27_y10),
    .I3(x28_y12)
);

(* keep, dont_touch *)
(* LOC = "X31/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110010000011)
) lut_31_7 (
    .O(x31_y7),
    .I0(x28_y10),
    .I1(x28_y6),
    .I2(1'b0),
    .I3(x29_y8)
);

(* keep, dont_touch *)
(* LOC = "X32/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000001010111)
) lut_32_7 (
    .O(x32_y7),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x29_y5),
    .I3(x30_y4)
);

(* keep, dont_touch *)
(* LOC = "X33/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000111111000)
) lut_33_7 (
    .O(x33_y7),
    .I0(x31_y5),
    .I1(x30_y9),
    .I2(x31_y9),
    .I3(x30_y12)
);

(* keep, dont_touch *)
(* LOC = "X34/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101110101001)
) lut_34_7 (
    .O(x34_y7),
    .I0(x32_y3),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X35/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010001010111)
) lut_35_7 (
    .O(x35_y7),
    .I0(1'b0),
    .I1(x33_y4),
    .I2(x32_y7),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X36/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111111010001)
) lut_36_7 (
    .O(x36_y7),
    .I0(x33_y5),
    .I1(x33_y6),
    .I2(x33_y8),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X37/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100110101110)
) lut_37_7 (
    .O(x37_y7),
    .I0(x34_y8),
    .I1(x35_y2),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X38/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111000011011)
) lut_38_7 (
    .O(x38_y7),
    .I0(x36_y4),
    .I1(x36_y7),
    .I2(x35_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X39/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011010100000)
) lut_39_7 (
    .O(x39_y7),
    .I0(x36_y5),
    .I1(1'b0),
    .I2(x36_y6),
    .I3(x37_y8)
);

(* keep, dont_touch *)
(* LOC = "X40/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111111010000)
) lut_40_7 (
    .O(x40_y7),
    .I0(x37_y6),
    .I1(1'b0),
    .I2(x38_y8),
    .I3(x38_y3)
);

(* keep, dont_touch *)
(* LOC = "X41/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100011011001)
) lut_41_7 (
    .O(x41_y7),
    .I0(1'b0),
    .I1(x38_y7),
    .I2(x39_y9),
    .I3(x38_y8)
);

(* keep, dont_touch *)
(* LOC = "X42/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000011101010)
) lut_42_7 (
    .O(x42_y7),
    .I0(1'b0),
    .I1(x40_y10),
    .I2(x39_y4),
    .I3(x39_y7)
);

(* keep, dont_touch *)
(* LOC = "X43/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001111110101)
) lut_43_7 (
    .O(x43_y7),
    .I0(x41_y4),
    .I1(x40_y4),
    .I2(x40_y3),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X44/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011100000010)
) lut_44_7 (
    .O(x44_y7),
    .I0(x41_y7),
    .I1(x41_y8),
    .I2(x41_y6),
    .I3(x42_y10)
);

(* keep, dont_touch *)
(* LOC = "X45/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101011011001)
) lut_45_7 (
    .O(x45_y7),
    .I0(x42_y12),
    .I1(x42_y6),
    .I2(x42_y10),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X46/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111001011001)
) lut_46_7 (
    .O(x46_y7),
    .I0(1'b0),
    .I1(x43_y5),
    .I2(x44_y10),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X47/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100000001100)
) lut_47_7 (
    .O(x47_y7),
    .I0(1'b0),
    .I1(x44_y5),
    .I2(x45_y5),
    .I3(x44_y4)
);

(* keep, dont_touch *)
(* LOC = "X48/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011001110110)
) lut_48_7 (
    .O(x48_y7),
    .I0(1'b0),
    .I1(x46_y12),
    .I2(x45_y3),
    .I3(x45_y11)
);

(* keep, dont_touch *)
(* LOC = "X49/Y7" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001010110011)
) lut_49_7 (
    .O(x49_y7),
    .I0(x46_y4),
    .I1(1'b0),
    .I2(x47_y6),
    .I3(x46_y6)
);

(* keep, dont_touch *)
(* LOC = "X0/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001001111011)
) lut_0_8 (
    .O(x0_y8),
    .I0(in9),
    .I1(1'b0),
    .I2(1'b0),
    .I3(in2)
);

(* keep, dont_touch *)
(* LOC = "X1/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100011110111)
) lut_1_8 (
    .O(x1_y8),
    .I0(1'b0),
    .I1(in1),
    .I2(in3),
    .I3(in9)
);

(* keep, dont_touch *)
(* LOC = "X2/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101000011000)
) lut_2_8 (
    .O(x2_y8),
    .I0(in3),
    .I1(in9),
    .I2(1'b0),
    .I3(in1)
);

(* keep, dont_touch *)
(* LOC = "X3/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101100100011)
) lut_3_8 (
    .O(x3_y8),
    .I0(x1_y3),
    .I1(1'b0),
    .I2(in7),
    .I3(in3)
);

(* keep, dont_touch *)
(* LOC = "X4/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101110111000)
) lut_4_8 (
    .O(x4_y8),
    .I0(x1_y12),
    .I1(x2_y9),
    .I2(x1_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X5/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000001111000)
) lut_5_8 (
    .O(x5_y8),
    .I0(1'b0),
    .I1(x3_y8),
    .I2(1'b0),
    .I3(x2_y10)
);

(* keep, dont_touch *)
(* LOC = "X6/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100110111110)
) lut_6_8 (
    .O(x6_y8),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x4_y12),
    .I3(x3_y4)
);

(* keep, dont_touch *)
(* LOC = "X7/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000000000100)
) lut_7_8 (
    .O(x7_y8),
    .I0(x5_y5),
    .I1(x5_y8),
    .I2(x5_y12),
    .I3(x5_y7)
);

(* keep, dont_touch *)
(* LOC = "X8/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000001011111)
) lut_8_8 (
    .O(x8_y8),
    .I0(x6_y10),
    .I1(x5_y7),
    .I2(x6_y7),
    .I3(x5_y3)
);

(* keep, dont_touch *)
(* LOC = "X9/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101110111110)
) lut_9_8 (
    .O(x9_y8),
    .I0(x6_y10),
    .I1(x6_y6),
    .I2(x6_y7),
    .I3(x5_y3)
);

(* keep, dont_touch *)
(* LOC = "X10/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000110111011)
) lut_10_8 (
    .O(x10_y8),
    .I0(x8_y11),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x7_y7)
);

(* keep, dont_touch *)
(* LOC = "X11/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110111111011)
) lut_11_8 (
    .O(x11_y8),
    .I0(1'b0),
    .I1(x8_y11),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X12/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001101011011)
) lut_12_8 (
    .O(x12_y8),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x10_y4),
    .I3(x9_y5)
);

(* keep, dont_touch *)
(* LOC = "X13/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001000001000)
) lut_13_8 (
    .O(x13_y8),
    .I0(x10_y8),
    .I1(x10_y6),
    .I2(1'b0),
    .I3(x11_y3)
);

(* keep, dont_touch *)
(* LOC = "X14/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010010111011)
) lut_14_8 (
    .O(x14_y8),
    .I0(x12_y7),
    .I1(x11_y13),
    .I2(x12_y7),
    .I3(x11_y12)
);

(* keep, dont_touch *)
(* LOC = "X15/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001011000110)
) lut_15_8 (
    .O(x15_y8),
    .I0(x12_y12),
    .I1(x13_y6),
    .I2(1'b0),
    .I3(x13_y5)
);

(* keep, dont_touch *)
(* LOC = "X16/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101111101000)
) lut_16_8 (
    .O(x16_y8),
    .I0(x14_y8),
    .I1(1'b0),
    .I2(x13_y3),
    .I3(x13_y7)
);

(* keep, dont_touch *)
(* LOC = "X17/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000101110111)
) lut_17_8 (
    .O(x17_y8),
    .I0(x15_y11),
    .I1(x15_y8),
    .I2(x15_y9),
    .I3(x15_y4)
);

(* keep, dont_touch *)
(* LOC = "X18/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100101001101)
) lut_18_8 (
    .O(x18_y8),
    .I0(x15_y5),
    .I1(x15_y9),
    .I2(x16_y8),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X19/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111000001110)
) lut_19_8 (
    .O(x19_y8),
    .I0(x17_y3),
    .I1(x17_y6),
    .I2(x16_y4),
    .I3(x16_y12)
);

(* keep, dont_touch *)
(* LOC = "X20/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110000000001)
) lut_20_8 (
    .O(x20_y8),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x18_y11)
);

(* keep, dont_touch *)
(* LOC = "X21/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010000011110)
) lut_21_8 (
    .O(x21_y8),
    .I0(x19_y6),
    .I1(x18_y4),
    .I2(x18_y10),
    .I3(x18_y3)
);

(* keep, dont_touch *)
(* LOC = "X22/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110110000101)
) lut_22_8 (
    .O(x22_y8),
    .I0(x20_y10),
    .I1(x19_y6),
    .I2(1'b0),
    .I3(x19_y10)
);

(* keep, dont_touch *)
(* LOC = "X23/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010011111100)
) lut_23_8 (
    .O(x23_y8),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x20_y12)
);

(* keep, dont_touch *)
(* LOC = "X24/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101111000001)
) lut_24_8 (
    .O(x24_y8),
    .I0(x21_y7),
    .I1(x22_y5),
    .I2(x22_y6),
    .I3(x21_y8)
);

(* keep, dont_touch *)
(* LOC = "X25/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111111101010)
) lut_25_8 (
    .O(x25_y8),
    .I0(x23_y12),
    .I1(x23_y3),
    .I2(1'b0),
    .I3(x23_y7)
);

(* keep, dont_touch *)
(* LOC = "X26/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001011100000)
) lut_26_8 (
    .O(x26_y8),
    .I0(x23_y13),
    .I1(x24_y6),
    .I2(x23_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X27/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001001111100)
) lut_27_8 (
    .O(x27_y8),
    .I0(x24_y8),
    .I1(x25_y7),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X28/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011100011010)
) lut_28_8 (
    .O(x28_y8),
    .I0(x26_y10),
    .I1(1'b0),
    .I2(x26_y10),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X29/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000100001110)
) lut_29_8 (
    .O(x29_y8),
    .I0(x27_y8),
    .I1(x26_y11),
    .I2(x27_y9),
    .I3(x27_y8)
);

(* keep, dont_touch *)
(* LOC = "X30/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001001111001)
) lut_30_8 (
    .O(x30_y8),
    .I0(x27_y11),
    .I1(x28_y8),
    .I2(x28_y13),
    .I3(x27_y9)
);

(* keep, dont_touch *)
(* LOC = "X31/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010101111000)
) lut_31_8 (
    .O(x31_y8),
    .I0(x28_y10),
    .I1(x29_y12),
    .I2(1'b0),
    .I3(x28_y11)
);

(* keep, dont_touch *)
(* LOC = "X32/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110100000101)
) lut_32_8 (
    .O(x32_y8),
    .I0(x29_y13),
    .I1(x29_y12),
    .I2(1'b0),
    .I3(x30_y4)
);

(* keep, dont_touch *)
(* LOC = "X33/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101111110011)
) lut_33_8 (
    .O(x33_y8),
    .I0(x31_y10),
    .I1(x30_y8),
    .I2(x31_y9),
    .I3(x31_y6)
);

(* keep, dont_touch *)
(* LOC = "X34/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100001101000)
) lut_34_8 (
    .O(x34_y8),
    .I0(x31_y10),
    .I1(x31_y13),
    .I2(x31_y7),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X35/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011111000010)
) lut_35_8 (
    .O(x35_y8),
    .I0(x32_y4),
    .I1(1'b0),
    .I2(x32_y9),
    .I3(x33_y12)
);

(* keep, dont_touch *)
(* LOC = "X36/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101011011001)
) lut_36_8 (
    .O(x36_y8),
    .I0(x34_y7),
    .I1(x33_y10),
    .I2(x33_y7),
    .I3(x33_y6)
);

(* keep, dont_touch *)
(* LOC = "X37/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100101110111)
) lut_37_8 (
    .O(x37_y8),
    .I0(x35_y9),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x34_y10)
);

(* keep, dont_touch *)
(* LOC = "X38/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000110110010)
) lut_38_8 (
    .O(x38_y8),
    .I0(x36_y8),
    .I1(x35_y12),
    .I2(x35_y9),
    .I3(x36_y3)
);

(* keep, dont_touch *)
(* LOC = "X39/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111100011111)
) lut_39_8 (
    .O(x39_y8),
    .I0(x37_y7),
    .I1(x37_y8),
    .I2(x36_y11),
    .I3(x37_y12)
);

(* keep, dont_touch *)
(* LOC = "X40/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111100101010)
) lut_40_8 (
    .O(x40_y8),
    .I0(x38_y13),
    .I1(x37_y3),
    .I2(x38_y9),
    .I3(x38_y13)
);

(* keep, dont_touch *)
(* LOC = "X41/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110110100001)
) lut_41_8 (
    .O(x41_y8),
    .I0(x39_y6),
    .I1(x38_y10),
    .I2(x38_y12),
    .I3(x39_y6)
);

(* keep, dont_touch *)
(* LOC = "X42/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001000111101)
) lut_42_8 (
    .O(x42_y8),
    .I0(x39_y8),
    .I1(x39_y8),
    .I2(x39_y3),
    .I3(x40_y7)
);

(* keep, dont_touch *)
(* LOC = "X43/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100100100111)
) lut_43_8 (
    .O(x43_y8),
    .I0(x41_y4),
    .I1(x41_y7),
    .I2(1'b0),
    .I3(x41_y11)
);

(* keep, dont_touch *)
(* LOC = "X44/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011000101101)
) lut_44_8 (
    .O(x44_y8),
    .I0(x41_y11),
    .I1(x41_y4),
    .I2(x42_y12),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X45/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000110010110)
) lut_45_8 (
    .O(x45_y8),
    .I0(x43_y5),
    .I1(x43_y4),
    .I2(x42_y11),
    .I3(x43_y7)
);

(* keep, dont_touch *)
(* LOC = "X46/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001100101011)
) lut_46_8 (
    .O(x46_y8),
    .I0(x43_y9),
    .I1(x43_y9),
    .I2(x44_y5),
    .I3(x43_y7)
);

(* keep, dont_touch *)
(* LOC = "X47/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100000110000)
) lut_47_8 (
    .O(x47_y8),
    .I0(x44_y5),
    .I1(x45_y8),
    .I2(x45_y4),
    .I3(x45_y4)
);

(* keep, dont_touch *)
(* LOC = "X48/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111101000110)
) lut_48_8 (
    .O(x48_y8),
    .I0(x45_y4),
    .I1(1'b0),
    .I2(x46_y10),
    .I3(x46_y12)
);

(* keep, dont_touch *)
(* LOC = "X49/Y8" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010110001000)
) lut_49_8 (
    .O(x49_y8),
    .I0(x46_y10),
    .I1(x46_y8),
    .I2(x47_y5),
    .I3(x46_y4)
);

(* keep, dont_touch *)
(* LOC = "X0/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101011111010)
) lut_0_9 (
    .O(x0_y9),
    .I0(1'b0),
    .I1(in9),
    .I2(in6),
    .I3(in6)
);

(* keep, dont_touch *)
(* LOC = "X1/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110011101011)
) lut_1_9 (
    .O(x1_y9),
    .I0(in8),
    .I1(1'b0),
    .I2(1'b0),
    .I3(in6)
);

(* keep, dont_touch *)
(* LOC = "X2/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110101001001)
) lut_2_9 (
    .O(x2_y9),
    .I0(in4),
    .I1(1'b0),
    .I2(1'b0),
    .I3(in5)
);

(* keep, dont_touch *)
(* LOC = "X3/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010111111011)
) lut_3_9 (
    .O(x3_y9),
    .I0(in5),
    .I1(in7),
    .I2(x1_y4),
    .I3(in6)
);

(* keep, dont_touch *)
(* LOC = "X4/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000010001111)
) lut_4_9 (
    .O(x4_y9),
    .I0(1'b0),
    .I1(x2_y13),
    .I2(x1_y7),
    .I3(x1_y8)
);

(* keep, dont_touch *)
(* LOC = "X5/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000000111110)
) lut_5_9 (
    .O(x5_y9),
    .I0(x3_y5),
    .I1(x2_y14),
    .I2(1'b0),
    .I3(x2_y14)
);

(* keep, dont_touch *)
(* LOC = "X6/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110100001010)
) lut_6_9 (
    .O(x6_y9),
    .I0(1'b0),
    .I1(x3_y10),
    .I2(x3_y5),
    .I3(x4_y11)
);

(* keep, dont_touch *)
(* LOC = "X7/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111000001001)
) lut_7_9 (
    .O(x7_y9),
    .I0(x5_y11),
    .I1(x4_y9),
    .I2(x4_y14),
    .I3(x4_y14)
);

(* keep, dont_touch *)
(* LOC = "X8/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100001101000)
) lut_8_9 (
    .O(x8_y9),
    .I0(x5_y4),
    .I1(x6_y7),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X9/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001101101011)
) lut_9_9 (
    .O(x9_y9),
    .I0(1'b0),
    .I1(x6_y13),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X10/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000001100011)
) lut_10_9 (
    .O(x10_y9),
    .I0(x7_y5),
    .I1(x7_y12),
    .I2(x7_y9),
    .I3(x8_y12)
);

(* keep, dont_touch *)
(* LOC = "X11/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110101001001)
) lut_11_9 (
    .O(x11_y9),
    .I0(x9_y10),
    .I1(x9_y9),
    .I2(x8_y8),
    .I3(x8_y13)
);

(* keep, dont_touch *)
(* LOC = "X12/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000011000100)
) lut_12_9 (
    .O(x12_y9),
    .I0(x10_y8),
    .I1(x9_y12),
    .I2(x10_y14),
    .I3(x9_y12)
);

(* keep, dont_touch *)
(* LOC = "X13/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011011101101)
) lut_13_9 (
    .O(x13_y9),
    .I0(x11_y7),
    .I1(x10_y8),
    .I2(x10_y8),
    .I3(x10_y4)
);

(* keep, dont_touch *)
(* LOC = "X14/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101111011000)
) lut_14_9 (
    .O(x14_y9),
    .I0(x11_y7),
    .I1(x11_y9),
    .I2(x12_y13),
    .I3(x12_y12)
);

(* keep, dont_touch *)
(* LOC = "X15/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010010110011)
) lut_15_9 (
    .O(x15_y9),
    .I0(x13_y4),
    .I1(x12_y14),
    .I2(1'b0),
    .I3(x13_y8)
);

(* keep, dont_touch *)
(* LOC = "X16/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010100010010)
) lut_16_9 (
    .O(x16_y9),
    .I0(x14_y8),
    .I1(x14_y10),
    .I2(x13_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X17/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110100000111)
) lut_17_9 (
    .O(x17_y9),
    .I0(x15_y8),
    .I1(x15_y7),
    .I2(x15_y14),
    .I3(x14_y12)
);

(* keep, dont_touch *)
(* LOC = "X18/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010011011010)
) lut_18_9 (
    .O(x18_y9),
    .I0(x15_y9),
    .I1(x15_y5),
    .I2(x16_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X19/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001101111001)
) lut_19_9 (
    .O(x19_y9),
    .I0(x17_y4),
    .I1(x17_y4),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X20/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111101001101)
) lut_20_9 (
    .O(x20_y9),
    .I0(x17_y14),
    .I1(x18_y5),
    .I2(1'b0),
    .I3(x17_y4)
);

(* keep, dont_touch *)
(* LOC = "X21/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011100111001)
) lut_21_9 (
    .O(x21_y9),
    .I0(x18_y4),
    .I1(1'b0),
    .I2(x19_y11),
    .I3(x19_y5)
);

(* keep, dont_touch *)
(* LOC = "X22/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111010010000)
) lut_22_9 (
    .O(x22_y9),
    .I0(x19_y10),
    .I1(x19_y9),
    .I2(x19_y4),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X23/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001110100101)
) lut_23_9 (
    .O(x23_y9),
    .I0(x20_y14),
    .I1(x20_y11),
    .I2(x20_y6),
    .I3(x21_y9)
);

(* keep, dont_touch *)
(* LOC = "X24/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010000111000)
) lut_24_9 (
    .O(x24_y9),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x21_y10),
    .I3(x22_y5)
);

(* keep, dont_touch *)
(* LOC = "X25/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100110111100)
) lut_25_9 (
    .O(x25_y9),
    .I0(x23_y4),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X26/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110110110101)
) lut_26_9 (
    .O(x26_y9),
    .I0(x24_y12),
    .I1(x24_y6),
    .I2(1'b0),
    .I3(x24_y5)
);

(* keep, dont_touch *)
(* LOC = "X27/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010110111101)
) lut_27_9 (
    .O(x27_y9),
    .I0(x25_y7),
    .I1(x24_y9),
    .I2(1'b0),
    .I3(x24_y10)
);

(* keep, dont_touch *)
(* LOC = "X28/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001101010101)
) lut_28_9 (
    .O(x28_y9),
    .I0(x25_y6),
    .I1(x25_y8),
    .I2(x25_y13),
    .I3(x26_y12)
);

(* keep, dont_touch *)
(* LOC = "X29/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110010001010)
) lut_29_9 (
    .O(x29_y9),
    .I0(x27_y8),
    .I1(x26_y8),
    .I2(x27_y14),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X30/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010100111100)
) lut_30_9 (
    .O(x30_y9),
    .I0(x27_y5),
    .I1(x27_y13),
    .I2(x27_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X31/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000010100111)
) lut_31_9 (
    .O(x31_y9),
    .I0(x28_y6),
    .I1(x28_y14),
    .I2(x29_y10),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X32/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000111101001)
) lut_32_9 (
    .O(x32_y9),
    .I0(x29_y12),
    .I1(x30_y12),
    .I2(x30_y7),
    .I3(x30_y13)
);

(* keep, dont_touch *)
(* LOC = "X33/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011000010011)
) lut_33_9 (
    .O(x33_y9),
    .I0(1'b0),
    .I1(x30_y14),
    .I2(1'b0),
    .I3(x30_y9)
);

(* keep, dont_touch *)
(* LOC = "X34/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111111000110)
) lut_34_9 (
    .O(x34_y9),
    .I0(1'b0),
    .I1(x31_y13),
    .I2(x32_y7),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X35/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010001100001)
) lut_35_9 (
    .O(x35_y9),
    .I0(1'b0),
    .I1(x33_y14),
    .I2(1'b0),
    .I3(x32_y11)
);

(* keep, dont_touch *)
(* LOC = "X36/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001011110111)
) lut_36_9 (
    .O(x36_y9),
    .I0(x33_y7),
    .I1(x33_y4),
    .I2(x33_y7),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X37/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100010100100)
) lut_37_9 (
    .O(x37_y9),
    .I0(x34_y7),
    .I1(x35_y13),
    .I2(x34_y6),
    .I3(x34_y4)
);

(* keep, dont_touch *)
(* LOC = "X38/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000011110110)
) lut_38_9 (
    .O(x38_y9),
    .I0(x35_y10),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x35_y12)
);

(* keep, dont_touch *)
(* LOC = "X39/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100001111110)
) lut_39_9 (
    .O(x39_y9),
    .I0(1'b0),
    .I1(x36_y13),
    .I2(x36_y5),
    .I3(x37_y13)
);

(* keep, dont_touch *)
(* LOC = "X40/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001000011001)
) lut_40_9 (
    .O(x40_y9),
    .I0(x38_y14),
    .I1(x37_y13),
    .I2(x37_y6),
    .I3(x37_y8)
);

(* keep, dont_touch *)
(* LOC = "X41/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001010101000)
) lut_41_9 (
    .O(x41_y9),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x39_y14),
    .I3(x38_y11)
);

(* keep, dont_touch *)
(* LOC = "X42/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110110110011)
) lut_42_9 (
    .O(x42_y9),
    .I0(1'b0),
    .I1(x39_y9),
    .I2(x39_y9),
    .I3(x40_y12)
);

(* keep, dont_touch *)
(* LOC = "X43/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111101111000)
) lut_43_9 (
    .O(x43_y9),
    .I0(x41_y6),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X44/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111011011100)
) lut_44_9 (
    .O(x44_y9),
    .I0(x41_y9),
    .I1(x42_y11),
    .I2(1'b0),
    .I3(x41_y5)
);

(* keep, dont_touch *)
(* LOC = "X45/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011101101000)
) lut_45_9 (
    .O(x45_y9),
    .I0(x43_y10),
    .I1(x43_y14),
    .I2(1'b0),
    .I3(x42_y10)
);

(* keep, dont_touch *)
(* LOC = "X46/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111001101011)
) lut_46_9 (
    .O(x46_y9),
    .I0(x43_y10),
    .I1(x43_y9),
    .I2(x44_y14),
    .I3(x44_y12)
);

(* keep, dont_touch *)
(* LOC = "X47/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001011010001)
) lut_47_9 (
    .O(x47_y9),
    .I0(x45_y8),
    .I1(x44_y11),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X48/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100001111010)
) lut_48_9 (
    .O(x48_y9),
    .I0(1'b0),
    .I1(x45_y6),
    .I2(x46_y5),
    .I3(x46_y6)
);

(* keep, dont_touch *)
(* LOC = "X49/Y9" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111101101010)
) lut_49_9 (
    .O(x49_y9),
    .I0(1'b0),
    .I1(x47_y8),
    .I2(x47_y13),
    .I3(x47_y10)
);

(* keep, dont_touch *)
(* LOC = "X0/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001000000101)
) lut_0_10 (
    .O(x0_y10),
    .I0(in0),
    .I1(in1),
    .I2(in0),
    .I3(in2)
);

(* keep, dont_touch *)
(* LOC = "X1/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011110110100)
) lut_1_10 (
    .O(x1_y10),
    .I0(1'b0),
    .I1(in9),
    .I2(1'b0),
    .I3(in7)
);

(* keep, dont_touch *)
(* LOC = "X2/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110110011010)
) lut_2_10 (
    .O(x2_y10),
    .I0(in7),
    .I1(in8),
    .I2(1'b0),
    .I3(in0)
);

(* keep, dont_touch *)
(* LOC = "X3/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011010101011)
) lut_3_10 (
    .O(x3_y10),
    .I0(x1_y15),
    .I1(x1_y6),
    .I2(x1_y7),
    .I3(in3)
);

(* keep, dont_touch *)
(* LOC = "X4/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101111010000)
) lut_4_10 (
    .O(x4_y10),
    .I0(x2_y15),
    .I1(x2_y6),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X5/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000110111011)
) lut_5_10 (
    .O(x5_y10),
    .I0(x2_y7),
    .I1(1'b0),
    .I2(x3_y15),
    .I3(x3_y11)
);

(* keep, dont_touch *)
(* LOC = "X6/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101011011111)
) lut_6_10 (
    .O(x6_y10),
    .I0(x3_y9),
    .I1(x4_y9),
    .I2(x4_y8),
    .I3(x3_y14)
);

(* keep, dont_touch *)
(* LOC = "X7/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110100000001)
) lut_7_10 (
    .O(x7_y10),
    .I0(x4_y12),
    .I1(x4_y13),
    .I2(x4_y8),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X8/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110101011111)
) lut_8_10 (
    .O(x8_y10),
    .I0(x6_y14),
    .I1(1'b0),
    .I2(x6_y9),
    .I3(x5_y6)
);

(* keep, dont_touch *)
(* LOC = "X9/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010010001011)
) lut_9_10 (
    .O(x9_y10),
    .I0(1'b0),
    .I1(x7_y9),
    .I2(x6_y9),
    .I3(x5_y6)
);

(* keep, dont_touch *)
(* LOC = "X10/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101011001011)
) lut_10_10 (
    .O(x10_y10),
    .I0(x7_y7),
    .I1(1'b0),
    .I2(x8_y13),
    .I3(x8_y5)
);

(* keep, dont_touch *)
(* LOC = "X11/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011110001010)
) lut_11_10 (
    .O(x11_y10),
    .I0(x8_y14),
    .I1(x9_y14),
    .I2(x9_y14),
    .I3(x8_y15)
);

(* keep, dont_touch *)
(* LOC = "X12/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010010011010)
) lut_12_10 (
    .O(x12_y10),
    .I0(x10_y7),
    .I1(x10_y5),
    .I2(1'b0),
    .I3(x9_y5)
);

(* keep, dont_touch *)
(* LOC = "X13/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110001110100)
) lut_13_10 (
    .O(x13_y10),
    .I0(x10_y8),
    .I1(x10_y7),
    .I2(1'b0),
    .I3(x10_y13)
);

(* keep, dont_touch *)
(* LOC = "X14/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100010000000)
) lut_14_10 (
    .O(x14_y10),
    .I0(x11_y14),
    .I1(x12_y9),
    .I2(x11_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X15/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010001111001)
) lut_15_10 (
    .O(x15_y10),
    .I0(x12_y11),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x12_y5)
);

(* keep, dont_touch *)
(* LOC = "X16/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000100111000)
) lut_16_10 (
    .O(x16_y10),
    .I0(x14_y14),
    .I1(x13_y14),
    .I2(x14_y11),
    .I3(x13_y9)
);

(* keep, dont_touch *)
(* LOC = "X17/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001000000010)
) lut_17_10 (
    .O(x17_y10),
    .I0(x15_y5),
    .I1(x14_y12),
    .I2(x14_y9),
    .I3(x14_y9)
);

(* keep, dont_touch *)
(* LOC = "X18/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001011101011)
) lut_18_10 (
    .O(x18_y10),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x16_y9),
    .I3(x15_y9)
);

(* keep, dont_touch *)
(* LOC = "X19/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001110111100)
) lut_19_10 (
    .O(x19_y10),
    .I0(x17_y7),
    .I1(1'b0),
    .I2(x16_y9),
    .I3(x17_y6)
);

(* keep, dont_touch *)
(* LOC = "X20/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011110000110)
) lut_20_10 (
    .O(x20_y10),
    .I0(x18_y10),
    .I1(x18_y10),
    .I2(x17_y7),
    .I3(x17_y10)
);

(* keep, dont_touch *)
(* LOC = "X21/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110000110000)
) lut_21_10 (
    .O(x21_y10),
    .I0(x19_y14),
    .I1(1'b0),
    .I2(x19_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X22/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111010001001)
) lut_22_10 (
    .O(x22_y10),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x20_y15),
    .I3(x19_y13)
);

(* keep, dont_touch *)
(* LOC = "X23/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001011111001)
) lut_23_10 (
    .O(x23_y10),
    .I0(1'b0),
    .I1(x21_y9),
    .I2(x21_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X24/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110100101101)
) lut_24_10 (
    .O(x24_y10),
    .I0(x21_y9),
    .I1(1'b0),
    .I2(x22_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X25/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001000010100)
) lut_25_10 (
    .O(x25_y10),
    .I0(x22_y13),
    .I1(x23_y5),
    .I2(x22_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X26/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101100010010)
) lut_26_10 (
    .O(x26_y10),
    .I0(x24_y12),
    .I1(x23_y14),
    .I2(x24_y15),
    .I3(x23_y13)
);

(* keep, dont_touch *)
(* LOC = "X27/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101100101101)
) lut_27_10 (
    .O(x27_y10),
    .I0(x24_y13),
    .I1(x25_y11),
    .I2(x25_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X28/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111011110100)
) lut_28_10 (
    .O(x28_y10),
    .I0(1'b0),
    .I1(x26_y9),
    .I2(x26_y8),
    .I3(x25_y14)
);

(* keep, dont_touch *)
(* LOC = "X29/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111110010101)
) lut_29_10 (
    .O(x29_y10),
    .I0(1'b0),
    .I1(x26_y7),
    .I2(x27_y7),
    .I3(x27_y10)
);

(* keep, dont_touch *)
(* LOC = "X30/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010100101001)
) lut_30_10 (
    .O(x30_y10),
    .I0(x28_y10),
    .I1(1'b0),
    .I2(x28_y13),
    .I3(x28_y15)
);

(* keep, dont_touch *)
(* LOC = "X31/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011101101110)
) lut_31_10 (
    .O(x31_y10),
    .I0(x29_y13),
    .I1(x29_y10),
    .I2(x29_y11),
    .I3(x28_y15)
);

(* keep, dont_touch *)
(* LOC = "X32/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110111101000)
) lut_32_10 (
    .O(x32_y10),
    .I0(x30_y9),
    .I1(1'b0),
    .I2(x29_y5),
    .I3(x29_y11)
);

(* keep, dont_touch *)
(* LOC = "X33/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111010011010)
) lut_33_10 (
    .O(x33_y10),
    .I0(x30_y6),
    .I1(x31_y9),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X34/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110011101100)
) lut_34_10 (
    .O(x34_y10),
    .I0(1'b0),
    .I1(x31_y9),
    .I2(x32_y5),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X35/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001101101011)
) lut_35_10 (
    .O(x35_y10),
    .I0(x32_y6),
    .I1(x32_y6),
    .I2(x32_y12),
    .I3(x33_y15)
);

(* keep, dont_touch *)
(* LOC = "X36/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101011100011)
) lut_36_10 (
    .O(x36_y10),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x33_y9),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X37/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000111101001)
) lut_37_10 (
    .O(x37_y10),
    .I0(x35_y12),
    .I1(x34_y5),
    .I2(1'b0),
    .I3(x35_y13)
);

(* keep, dont_touch *)
(* LOC = "X38/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001100101001)
) lut_38_10 (
    .O(x38_y10),
    .I0(x35_y7),
    .I1(x36_y14),
    .I2(x35_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X39/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011100100110)
) lut_39_10 (
    .O(x39_y10),
    .I0(x36_y7),
    .I1(x36_y14),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X40/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111101111000)
) lut_40_10 (
    .O(x40_y10),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x38_y11),
    .I3(x38_y7)
);

(* keep, dont_touch *)
(* LOC = "X41/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011001011010)
) lut_41_10 (
    .O(x41_y10),
    .I0(x39_y15),
    .I1(x38_y10),
    .I2(x38_y5),
    .I3(x38_y13)
);

(* keep, dont_touch *)
(* LOC = "X42/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011011101000)
) lut_42_10 (
    .O(x42_y10),
    .I0(x39_y11),
    .I1(x40_y10),
    .I2(x40_y9),
    .I3(x40_y9)
);

(* keep, dont_touch *)
(* LOC = "X43/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110111010010)
) lut_43_10 (
    .O(x43_y10),
    .I0(x40_y15),
    .I1(x41_y11),
    .I2(x41_y10),
    .I3(x41_y9)
);

(* keep, dont_touch *)
(* LOC = "X44/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011000100101)
) lut_44_10 (
    .O(x44_y10),
    .I0(x42_y15),
    .I1(x42_y12),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X45/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011010000000)
) lut_45_10 (
    .O(x45_y10),
    .I0(x42_y7),
    .I1(x42_y9),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X46/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001011100101)
) lut_46_10 (
    .O(x46_y10),
    .I0(1'b0),
    .I1(x43_y14),
    .I2(x43_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X47/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100111101111)
) lut_47_10 (
    .O(x47_y10),
    .I0(x45_y14),
    .I1(1'b0),
    .I2(x44_y8),
    .I3(x44_y6)
);

(* keep, dont_touch *)
(* LOC = "X48/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101110011100)
) lut_48_10 (
    .O(x48_y10),
    .I0(1'b0),
    .I1(x46_y14),
    .I2(x45_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X49/Y10" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111101110011)
) lut_49_10 (
    .O(x49_y10),
    .I0(x46_y11),
    .I1(x47_y13),
    .I2(1'b0),
    .I3(x47_y14)
);

(* keep, dont_touch *)
(* LOC = "X0/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111111010100)
) lut_0_11 (
    .O(x0_y11),
    .I0(in6),
    .I1(in7),
    .I2(1'b0),
    .I3(in7)
);

(* keep, dont_touch *)
(* LOC = "X1/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011110100110)
) lut_1_11 (
    .O(x1_y11),
    .I0(in9),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X2/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110110100011)
) lut_2_11 (
    .O(x2_y11),
    .I0(in8),
    .I1(1'b0),
    .I2(in6),
    .I3(in6)
);

(* keep, dont_touch *)
(* LOC = "X3/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000010000010)
) lut_3_11 (
    .O(x3_y11),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(in2)
);

(* keep, dont_touch *)
(* LOC = "X4/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110110101000)
) lut_4_11 (
    .O(x4_y11),
    .I0(x1_y8),
    .I1(x2_y8),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X5/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100111010010)
) lut_5_11 (
    .O(x5_y11),
    .I0(x3_y10),
    .I1(1'b0),
    .I2(x2_y9),
    .I3(x3_y16)
);

(* keep, dont_touch *)
(* LOC = "X6/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100101100010)
) lut_6_11 (
    .O(x6_y11),
    .I0(x4_y15),
    .I1(x3_y16),
    .I2(x4_y14),
    .I3(x4_y6)
);

(* keep, dont_touch *)
(* LOC = "X7/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110000111001)
) lut_7_11 (
    .O(x7_y11),
    .I0(x5_y8),
    .I1(x5_y7),
    .I2(1'b0),
    .I3(x5_y11)
);

(* keep, dont_touch *)
(* LOC = "X8/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010010110101)
) lut_8_11 (
    .O(x8_y11),
    .I0(x5_y8),
    .I1(x6_y9),
    .I2(x5_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X9/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100011110011)
) lut_9_11 (
    .O(x9_y11),
    .I0(x7_y8),
    .I1(x6_y16),
    .I2(x5_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X10/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011110000110)
) lut_10_11 (
    .O(x10_y11),
    .I0(1'b0),
    .I1(x8_y10),
    .I2(1'b0),
    .I3(x7_y15)
);

(* keep, dont_touch *)
(* LOC = "X11/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101100000000)
) lut_11_11 (
    .O(x11_y11),
    .I0(x9_y16),
    .I1(1'b0),
    .I2(x9_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X12/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011111001010)
) lut_12_11 (
    .O(x12_y11),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x10_y6),
    .I3(x10_y16)
);

(* keep, dont_touch *)
(* LOC = "X13/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101110010001)
) lut_13_11 (
    .O(x13_y11),
    .I0(x11_y14),
    .I1(1'b0),
    .I2(x10_y11),
    .I3(x10_y10)
);

(* keep, dont_touch *)
(* LOC = "X14/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011100000110)
) lut_14_11 (
    .O(x14_y11),
    .I0(x12_y8),
    .I1(x11_y11),
    .I2(x12_y8),
    .I3(x11_y15)
);

(* keep, dont_touch *)
(* LOC = "X15/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011000000001)
) lut_15_11 (
    .O(x15_y11),
    .I0(x12_y7),
    .I1(x13_y8),
    .I2(x12_y6),
    .I3(x12_y11)
);

(* keep, dont_touch *)
(* LOC = "X16/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110101111011)
) lut_16_11 (
    .O(x16_y11),
    .I0(x13_y11),
    .I1(x13_y8),
    .I2(x14_y10),
    .I3(x14_y16)
);

(* keep, dont_touch *)
(* LOC = "X17/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110001000100)
) lut_17_11 (
    .O(x17_y11),
    .I0(x15_y10),
    .I1(x15_y16),
    .I2(x15_y12),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X18/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100000110100)
) lut_18_11 (
    .O(x18_y11),
    .I0(1'b0),
    .I1(x16_y6),
    .I2(x15_y15),
    .I3(x15_y9)
);

(* keep, dont_touch *)
(* LOC = "X19/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111111000001)
) lut_19_11 (
    .O(x19_y11),
    .I0(x17_y14),
    .I1(x17_y8),
    .I2(x17_y11),
    .I3(x16_y8)
);

(* keep, dont_touch *)
(* LOC = "X20/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011010101000)
) lut_20_11 (
    .O(x20_y11),
    .I0(x17_y13),
    .I1(x17_y8),
    .I2(x17_y15),
    .I3(x18_y6)
);

(* keep, dont_touch *)
(* LOC = "X21/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100100111000)
) lut_21_11 (
    .O(x21_y11),
    .I0(1'b0),
    .I1(x19_y10),
    .I2(1'b0),
    .I3(x18_y14)
);

(* keep, dont_touch *)
(* LOC = "X22/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111011111000)
) lut_22_11 (
    .O(x22_y11),
    .I0(x19_y8),
    .I1(x19_y16),
    .I2(x19_y12),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X23/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100111101010)
) lut_23_11 (
    .O(x23_y11),
    .I0(x20_y11),
    .I1(x21_y9),
    .I2(x20_y6),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X24/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100001100000)
) lut_24_11 (
    .O(x24_y11),
    .I0(x21_y8),
    .I1(x22_y8),
    .I2(x22_y9),
    .I3(x21_y12)
);

(* keep, dont_touch *)
(* LOC = "X25/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000000001011)
) lut_25_11 (
    .O(x25_y11),
    .I0(x22_y6),
    .I1(x23_y15),
    .I2(x23_y10),
    .I3(x23_y10)
);

(* keep, dont_touch *)
(* LOC = "X26/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110010011110)
) lut_26_11 (
    .O(x26_y11),
    .I0(x23_y13),
    .I1(1'b0),
    .I2(x24_y12),
    .I3(x24_y16)
);

(* keep, dont_touch *)
(* LOC = "X27/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001011000001)
) lut_27_11 (
    .O(x27_y11),
    .I0(x24_y9),
    .I1(1'b0),
    .I2(x25_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X28/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100111101001)
) lut_28_11 (
    .O(x28_y11),
    .I0(1'b0),
    .I1(x26_y12),
    .I2(x25_y7),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X29/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100100110011)
) lut_29_11 (
    .O(x29_y11),
    .I0(1'b0),
    .I1(x26_y6),
    .I2(x27_y14),
    .I3(x27_y10)
);

(* keep, dont_touch *)
(* LOC = "X30/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011100110000)
) lut_30_11 (
    .O(x30_y11),
    .I0(1'b0),
    .I1(x27_y9),
    .I2(1'b0),
    .I3(x27_y9)
);

(* keep, dont_touch *)
(* LOC = "X31/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010111100000)
) lut_31_11 (
    .O(x31_y11),
    .I0(x28_y11),
    .I1(x29_y11),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X32/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001001001100)
) lut_32_11 (
    .O(x32_y11),
    .I0(1'b0),
    .I1(x29_y15),
    .I2(x30_y10),
    .I3(x30_y11)
);

(* keep, dont_touch *)
(* LOC = "X33/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000100111010)
) lut_33_11 (
    .O(x33_y11),
    .I0(x31_y9),
    .I1(x31_y13),
    .I2(x31_y8),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X34/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110110001100)
) lut_34_11 (
    .O(x34_y11),
    .I0(1'b0),
    .I1(x32_y6),
    .I2(x31_y12),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X35/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111001110000)
) lut_35_11 (
    .O(x35_y11),
    .I0(x32_y7),
    .I1(x32_y8),
    .I2(1'b0),
    .I3(x32_y13)
);

(* keep, dont_touch *)
(* LOC = "X36/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111100000001)
) lut_36_11 (
    .O(x36_y11),
    .I0(x34_y9),
    .I1(1'b0),
    .I2(x34_y10),
    .I3(x33_y10)
);

(* keep, dont_touch *)
(* LOC = "X37/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100001011101)
) lut_37_11 (
    .O(x37_y11),
    .I0(x35_y12),
    .I1(x34_y15),
    .I2(x35_y10),
    .I3(x35_y10)
);

(* keep, dont_touch *)
(* LOC = "X38/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010111010100)
) lut_38_11 (
    .O(x38_y11),
    .I0(x35_y11),
    .I1(x36_y9),
    .I2(1'b0),
    .I3(x35_y15)
);

(* keep, dont_touch *)
(* LOC = "X39/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101111010111)
) lut_39_11 (
    .O(x39_y11),
    .I0(x37_y13),
    .I1(1'b0),
    .I2(x36_y8),
    .I3(x37_y13)
);

(* keep, dont_touch *)
(* LOC = "X40/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001001110101)
) lut_40_11 (
    .O(x40_y11),
    .I0(x38_y16),
    .I1(x38_y15),
    .I2(1'b0),
    .I3(x38_y9)
);

(* keep, dont_touch *)
(* LOC = "X41/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100100001001)
) lut_41_11 (
    .O(x41_y11),
    .I0(x38_y10),
    .I1(x39_y10),
    .I2(x39_y9),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X42/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011110011111)
) lut_42_11 (
    .O(x42_y11),
    .I0(x40_y14),
    .I1(1'b0),
    .I2(x39_y10),
    .I3(x40_y15)
);

(* keep, dont_touch *)
(* LOC = "X43/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000010101100)
) lut_43_11 (
    .O(x43_y11),
    .I0(x41_y14),
    .I1(x41_y11),
    .I2(1'b0),
    .I3(x40_y7)
);

(* keep, dont_touch *)
(* LOC = "X44/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011000011001)
) lut_44_11 (
    .O(x44_y11),
    .I0(1'b0),
    .I1(x42_y11),
    .I2(x41_y6),
    .I3(x41_y13)
);

(* keep, dont_touch *)
(* LOC = "X45/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010010101001)
) lut_45_11 (
    .O(x45_y11),
    .I0(x43_y16),
    .I1(1'b0),
    .I2(x43_y12),
    .I3(x42_y13)
);

(* keep, dont_touch *)
(* LOC = "X46/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011010100000)
) lut_46_11 (
    .O(x46_y11),
    .I0(1'b0),
    .I1(x43_y16),
    .I2(1'b0),
    .I3(x43_y10)
);

(* keep, dont_touch *)
(* LOC = "X47/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011100011011)
) lut_47_11 (
    .O(x47_y11),
    .I0(x44_y13),
    .I1(x44_y15),
    .I2(x44_y14),
    .I3(x44_y9)
);

(* keep, dont_touch *)
(* LOC = "X48/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110100000100)
) lut_48_11 (
    .O(x48_y11),
    .I0(x46_y9),
    .I1(x46_y8),
    .I2(1'b0),
    .I3(x46_y16)
);

(* keep, dont_touch *)
(* LOC = "X49/Y11" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000000010100)
) lut_49_11 (
    .O(x49_y11),
    .I0(x46_y13),
    .I1(x46_y9),
    .I2(x46_y10),
    .I3(x46_y16)
);

(* keep, dont_touch *)
(* LOC = "X0/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101100001001)
) lut_0_12 (
    .O(x0_y12),
    .I0(in8),
    .I1(1'b0),
    .I2(1'b0),
    .I3(in2)
);

(* keep, dont_touch *)
(* LOC = "X1/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111000101100)
) lut_1_12 (
    .O(x1_y12),
    .I0(in4),
    .I1(in8),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X2/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100000101110)
) lut_2_12 (
    .O(x2_y12),
    .I0(in9),
    .I1(1'b0),
    .I2(in0),
    .I3(in2)
);

(* keep, dont_touch *)
(* LOC = "X3/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011111110100)
) lut_3_12 (
    .O(x3_y12),
    .I0(in6),
    .I1(1'b0),
    .I2(x1_y11),
    .I3(in6)
);

(* keep, dont_touch *)
(* LOC = "X4/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111100011001)
) lut_4_12 (
    .O(x4_y12),
    .I0(x1_y12),
    .I1(x2_y14),
    .I2(x2_y13),
    .I3(x2_y17)
);

(* keep, dont_touch *)
(* LOC = "X5/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110110100001)
) lut_5_12 (
    .O(x5_y12),
    .I0(x2_y17),
    .I1(x3_y8),
    .I2(x2_y14),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X6/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000101010010)
) lut_6_12 (
    .O(x6_y12),
    .I0(x4_y17),
    .I1(x3_y15),
    .I2(1'b0),
    .I3(x4_y11)
);

(* keep, dont_touch *)
(* LOC = "X7/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101110000100)
) lut_7_12 (
    .O(x7_y12),
    .I0(x4_y7),
    .I1(1'b0),
    .I2(x4_y8),
    .I3(x5_y10)
);

(* keep, dont_touch *)
(* LOC = "X8/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010001100010)
) lut_8_12 (
    .O(x8_y12),
    .I0(x6_y15),
    .I1(x5_y9),
    .I2(x5_y10),
    .I3(x5_y17)
);

(* keep, dont_touch *)
(* LOC = "X9/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000010110000)
) lut_9_12 (
    .O(x9_y12),
    .I0(x6_y16),
    .I1(x6_y10),
    .I2(x5_y10),
    .I3(x5_y17)
);

(* keep, dont_touch *)
(* LOC = "X10/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001010110011)
) lut_10_12 (
    .O(x10_y12),
    .I0(x7_y16),
    .I1(x7_y17),
    .I2(1'b0),
    .I3(x8_y9)
);

(* keep, dont_touch *)
(* LOC = "X11/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101110010110)
) lut_11_12 (
    .O(x11_y12),
    .I0(1'b0),
    .I1(x9_y9),
    .I2(x9_y14),
    .I3(x8_y17)
);

(* keep, dont_touch *)
(* LOC = "X12/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111100001001)
) lut_12_12 (
    .O(x12_y12),
    .I0(x9_y16),
    .I1(x9_y12),
    .I2(x9_y10),
    .I3(x9_y16)
);

(* keep, dont_touch *)
(* LOC = "X13/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010111100010)
) lut_13_12 (
    .O(x13_y12),
    .I0(x11_y17),
    .I1(x11_y13),
    .I2(x11_y13),
    .I3(x10_y13)
);

(* keep, dont_touch *)
(* LOC = "X14/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110010000000)
) lut_14_12 (
    .O(x14_y12),
    .I0(1'b0),
    .I1(x12_y8),
    .I2(x11_y11),
    .I3(x11_y17)
);

(* keep, dont_touch *)
(* LOC = "X15/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100101101101)
) lut_15_12 (
    .O(x15_y12),
    .I0(1'b0),
    .I1(x12_y12),
    .I2(x13_y16),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X16/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110011001011)
) lut_16_12 (
    .O(x16_y12),
    .I0(x14_y15),
    .I1(x14_y11),
    .I2(x14_y12),
    .I3(x13_y10)
);

(* keep, dont_touch *)
(* LOC = "X17/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111011110101)
) lut_17_12 (
    .O(x17_y12),
    .I0(x14_y9),
    .I1(x15_y8),
    .I2(1'b0),
    .I3(x14_y15)
);

(* keep, dont_touch *)
(* LOC = "X18/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001111001100)
) lut_18_12 (
    .O(x18_y12),
    .I0(1'b0),
    .I1(x15_y7),
    .I2(1'b0),
    .I3(x16_y7)
);

(* keep, dont_touch *)
(* LOC = "X19/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100001011011)
) lut_19_12 (
    .O(x19_y12),
    .I0(x16_y8),
    .I1(1'b0),
    .I2(x16_y8),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X20/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110100011101)
) lut_20_12 (
    .O(x20_y12),
    .I0(1'b0),
    .I1(x17_y14),
    .I2(x17_y10),
    .I3(x18_y12)
);

(* keep, dont_touch *)
(* LOC = "X21/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110001001000)
) lut_21_12 (
    .O(x21_y12),
    .I0(x18_y10),
    .I1(x19_y17),
    .I2(x18_y15),
    .I3(x18_y13)
);

(* keep, dont_touch *)
(* LOC = "X22/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100111101011)
) lut_22_12 (
    .O(x22_y12),
    .I0(x19_y9),
    .I1(x19_y12),
    .I2(x19_y17),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X23/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000001111111)
) lut_23_12 (
    .O(x23_y12),
    .I0(x21_y8),
    .I1(1'b0),
    .I2(x21_y14),
    .I3(x21_y11)
);

(* keep, dont_touch *)
(* LOC = "X24/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100010100101)
) lut_24_12 (
    .O(x24_y12),
    .I0(x22_y17),
    .I1(1'b0),
    .I2(x22_y16),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X25/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001011000111)
) lut_25_12 (
    .O(x25_y12),
    .I0(x22_y11),
    .I1(x22_y17),
    .I2(x23_y10),
    .I3(x22_y7)
);

(* keep, dont_touch *)
(* LOC = "X26/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111111110100)
) lut_26_12 (
    .O(x26_y12),
    .I0(x23_y7),
    .I1(1'b0),
    .I2(x23_y11),
    .I3(x24_y12)
);

(* keep, dont_touch *)
(* LOC = "X27/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011001011011)
) lut_27_12 (
    .O(x27_y12),
    .I0(x24_y15),
    .I1(x25_y17),
    .I2(x25_y16),
    .I3(x24_y11)
);

(* keep, dont_touch *)
(* LOC = "X28/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001101011000)
) lut_28_12 (
    .O(x28_y12),
    .I0(x26_y12),
    .I1(x26_y10),
    .I2(1'b0),
    .I3(x26_y9)
);

(* keep, dont_touch *)
(* LOC = "X29/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010000011110)
) lut_29_12 (
    .O(x29_y12),
    .I0(1'b0),
    .I1(x26_y8),
    .I2(x27_y8),
    .I3(x26_y13)
);

(* keep, dont_touch *)
(* LOC = "X30/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001110111100)
) lut_30_12 (
    .O(x30_y12),
    .I0(x27_y17),
    .I1(x28_y9),
    .I2(x27_y16),
    .I3(x28_y10)
);

(* keep, dont_touch *)
(* LOC = "X31/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010100101110)
) lut_31_12 (
    .O(x31_y12),
    .I0(1'b0),
    .I1(x28_y13),
    .I2(x28_y14),
    .I3(x28_y14)
);

(* keep, dont_touch *)
(* LOC = "X32/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000101111001)
) lut_32_12 (
    .O(x32_y12),
    .I0(1'b0),
    .I1(x29_y12),
    .I2(x29_y17),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X33/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101010100101)
) lut_33_12 (
    .O(x33_y12),
    .I0(x31_y7),
    .I1(x30_y9),
    .I2(x31_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X34/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101010010100)
) lut_34_12 (
    .O(x34_y12),
    .I0(x32_y14),
    .I1(1'b0),
    .I2(x32_y9),
    .I3(x31_y12)
);

(* keep, dont_touch *)
(* LOC = "X35/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100111000100)
) lut_35_12 (
    .O(x35_y12),
    .I0(1'b0),
    .I1(x33_y15),
    .I2(x33_y9),
    .I3(x33_y10)
);

(* keep, dont_touch *)
(* LOC = "X36/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111100101001)
) lut_36_12 (
    .O(x36_y12),
    .I0(x34_y7),
    .I1(x33_y8),
    .I2(x33_y7),
    .I3(x34_y15)
);

(* keep, dont_touch *)
(* LOC = "X37/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010010000110)
) lut_37_12 (
    .O(x37_y12),
    .I0(x34_y7),
    .I1(x34_y13),
    .I2(1'b0),
    .I3(x35_y9)
);

(* keep, dont_touch *)
(* LOC = "X38/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000111010101)
) lut_38_12 (
    .O(x38_y12),
    .I0(x35_y9),
    .I1(x36_y9),
    .I2(x35_y14),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X39/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111000011000)
) lut_39_12 (
    .O(x39_y12),
    .I0(x36_y14),
    .I1(1'b0),
    .I2(x37_y11),
    .I3(x37_y9)
);

(* keep, dont_touch *)
(* LOC = "X40/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000011000000)
) lut_40_12 (
    .O(x40_y12),
    .I0(1'b0),
    .I1(x37_y15),
    .I2(1'b0),
    .I3(x37_y7)
);

(* keep, dont_touch *)
(* LOC = "X41/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100000010100)
) lut_41_12 (
    .O(x41_y12),
    .I0(x39_y12),
    .I1(x39_y10),
    .I2(x38_y16),
    .I3(x39_y13)
);

(* keep, dont_touch *)
(* LOC = "X42/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101011111000)
) lut_42_12 (
    .O(x42_y12),
    .I0(x40_y10),
    .I1(1'b0),
    .I2(x40_y11),
    .I3(x39_y7)
);

(* keep, dont_touch *)
(* LOC = "X43/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011000111011)
) lut_43_12 (
    .O(x43_y12),
    .I0(x40_y17),
    .I1(x40_y14),
    .I2(x40_y14),
    .I3(x40_y9)
);

(* keep, dont_touch *)
(* LOC = "X44/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111001110100)
) lut_44_12 (
    .O(x44_y12),
    .I0(x41_y12),
    .I1(x41_y14),
    .I2(x42_y14),
    .I3(x41_y11)
);

(* keep, dont_touch *)
(* LOC = "X45/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011100110111)
) lut_45_12 (
    .O(x45_y12),
    .I0(x42_y17),
    .I1(1'b0),
    .I2(x42_y9),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X46/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001100110000)
) lut_46_12 (
    .O(x46_y12),
    .I0(1'b0),
    .I1(x44_y11),
    .I2(x44_y10),
    .I3(x44_y14)
);

(* keep, dont_touch *)
(* LOC = "X47/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001101010101)
) lut_47_12 (
    .O(x47_y12),
    .I0(x44_y8),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x44_y15)
);

(* keep, dont_touch *)
(* LOC = "X48/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110100101101)
) lut_48_12 (
    .O(x48_y12),
    .I0(x46_y10),
    .I1(x45_y16),
    .I2(x46_y15),
    .I3(x45_y15)
);

(* keep, dont_touch *)
(* LOC = "X49/Y12" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101111111111)
) lut_49_12 (
    .O(x49_y12),
    .I0(x47_y9),
    .I1(x47_y7),
    .I2(1'b0),
    .I3(x47_y7)
);

(* keep, dont_touch *)
(* LOC = "X0/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001100011001)
) lut_0_13 (
    .O(x0_y13),
    .I0(1'b0),
    .I1(in2),
    .I2(in2),
    .I3(in7)
);

(* keep, dont_touch *)
(* LOC = "X1/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000011000100)
) lut_1_13 (
    .O(x1_y13),
    .I0(in7),
    .I1(1'b0),
    .I2(1'b0),
    .I3(in1)
);

(* keep, dont_touch *)
(* LOC = "X2/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010010101100)
) lut_2_13 (
    .O(x2_y13),
    .I0(in4),
    .I1(in3),
    .I2(in2),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X3/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011001101011)
) lut_3_13 (
    .O(x3_y13),
    .I0(x1_y18),
    .I1(x1_y9),
    .I2(x1_y13),
    .I3(in5)
);

(* keep, dont_touch *)
(* LOC = "X4/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110001100101)
) lut_4_13 (
    .O(x4_y13),
    .I0(x2_y9),
    .I1(1'b0),
    .I2(x2_y10),
    .I3(x1_y14)
);

(* keep, dont_touch *)
(* LOC = "X5/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100111010111)
) lut_5_13 (
    .O(x5_y13),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x3_y16),
    .I3(x2_y18)
);

(* keep, dont_touch *)
(* LOC = "X6/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101011001000)
) lut_6_13 (
    .O(x6_y13),
    .I0(x3_y11),
    .I1(x3_y8),
    .I2(x4_y9),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X7/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100010000100)
) lut_7_13 (
    .O(x7_y13),
    .I0(x5_y17),
    .I1(x5_y17),
    .I2(x5_y9),
    .I3(x4_y12)
);

(* keep, dont_touch *)
(* LOC = "X8/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110011010111)
) lut_8_13 (
    .O(x8_y13),
    .I0(x5_y13),
    .I1(1'b0),
    .I2(x6_y13),
    .I3(x6_y15)
);

(* keep, dont_touch *)
(* LOC = "X9/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010000001100)
) lut_9_13 (
    .O(x9_y13),
    .I0(1'b0),
    .I1(x6_y8),
    .I2(x6_y13),
    .I3(x6_y15)
);

(* keep, dont_touch *)
(* LOC = "X10/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100000110011)
) lut_10_13 (
    .O(x10_y13),
    .I0(x8_y13),
    .I1(1'b0),
    .I2(x8_y10),
    .I3(x7_y12)
);

(* keep, dont_touch *)
(* LOC = "X11/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001000111000)
) lut_11_13 (
    .O(x11_y13),
    .I0(1'b0),
    .I1(x9_y11),
    .I2(x8_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X12/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111100110100)
) lut_12_13 (
    .O(x12_y13),
    .I0(x10_y10),
    .I1(x10_y16),
    .I2(x9_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X13/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000010011011)
) lut_13_13 (
    .O(x13_y13),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x10_y18),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X14/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111111101111)
) lut_14_13 (
    .O(x14_y13),
    .I0(1'b0),
    .I1(x12_y15),
    .I2(x11_y16),
    .I3(x12_y18)
);

(* keep, dont_touch *)
(* LOC = "X15/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110101100011)
) lut_15_13 (
    .O(x15_y13),
    .I0(x12_y17),
    .I1(x12_y9),
    .I2(x12_y13),
    .I3(x13_y10)
);

(* keep, dont_touch *)
(* LOC = "X16/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110001101011)
) lut_16_13 (
    .O(x16_y13),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x13_y13),
    .I3(x14_y15)
);

(* keep, dont_touch *)
(* LOC = "X17/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010101000001)
) lut_17_13 (
    .O(x17_y13),
    .I0(x14_y12),
    .I1(x14_y11),
    .I2(x14_y16),
    .I3(x14_y15)
);

(* keep, dont_touch *)
(* LOC = "X18/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100011010101)
) lut_18_13 (
    .O(x18_y13),
    .I0(x16_y14),
    .I1(x16_y9),
    .I2(x16_y17),
    .I3(x15_y8)
);

(* keep, dont_touch *)
(* LOC = "X19/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100110100011)
) lut_19_13 (
    .O(x19_y13),
    .I0(x16_y13),
    .I1(1'b0),
    .I2(x16_y10),
    .I3(x16_y16)
);

(* keep, dont_touch *)
(* LOC = "X20/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011101101100)
) lut_20_13 (
    .O(x20_y13),
    .I0(1'b0),
    .I1(x18_y14),
    .I2(x17_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X21/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011011101111)
) lut_21_13 (
    .O(x21_y13),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x19_y8),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X22/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000010100100)
) lut_22_13 (
    .O(x22_y13),
    .I0(x19_y9),
    .I1(x20_y8),
    .I2(x20_y9),
    .I3(x19_y18)
);

(* keep, dont_touch *)
(* LOC = "X23/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100010010010)
) lut_23_13 (
    .O(x23_y13),
    .I0(1'b0),
    .I1(x21_y16),
    .I2(x21_y12),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X24/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100000111011)
) lut_24_13 (
    .O(x24_y13),
    .I0(x22_y12),
    .I1(x21_y8),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X25/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000111110010)
) lut_25_13 (
    .O(x25_y13),
    .I0(1'b0),
    .I1(x23_y10),
    .I2(x22_y12),
    .I3(x23_y15)
);

(* keep, dont_touch *)
(* LOC = "X26/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010000001100)
) lut_26_13 (
    .O(x26_y13),
    .I0(1'b0),
    .I1(x23_y12),
    .I2(x23_y12),
    .I3(x24_y8)
);

(* keep, dont_touch *)
(* LOC = "X27/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001011100111)
) lut_27_13 (
    .O(x27_y13),
    .I0(x25_y16),
    .I1(x24_y10),
    .I2(x25_y11),
    .I3(x24_y14)
);

(* keep, dont_touch *)
(* LOC = "X28/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001001011111)
) lut_28_13 (
    .O(x28_y13),
    .I0(x25_y11),
    .I1(1'b0),
    .I2(x26_y10),
    .I3(x26_y15)
);

(* keep, dont_touch *)
(* LOC = "X29/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011100110010)
) lut_29_13 (
    .O(x29_y13),
    .I0(x27_y11),
    .I1(x27_y14),
    .I2(x27_y17),
    .I3(x27_y17)
);

(* keep, dont_touch *)
(* LOC = "X30/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001111100100)
) lut_30_13 (
    .O(x30_y13),
    .I0(x28_y9),
    .I1(x28_y12),
    .I2(x27_y17),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X31/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110101101000)
) lut_31_13 (
    .O(x31_y13),
    .I0(x28_y8),
    .I1(1'b0),
    .I2(x28_y17),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X32/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101001110000)
) lut_32_13 (
    .O(x32_y13),
    .I0(x30_y13),
    .I1(x30_y14),
    .I2(x30_y14),
    .I3(x29_y9)
);

(* keep, dont_touch *)
(* LOC = "X33/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100101000101)
) lut_33_13 (
    .O(x33_y13),
    .I0(x31_y8),
    .I1(x30_y15),
    .I2(x30_y10),
    .I3(x31_y11)
);

(* keep, dont_touch *)
(* LOC = "X34/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101010110110)
) lut_34_13 (
    .O(x34_y13),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x32_y8)
);

(* keep, dont_touch *)
(* LOC = "X35/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000001010110)
) lut_35_13 (
    .O(x35_y13),
    .I0(x33_y8),
    .I1(x33_y18),
    .I2(x32_y17),
    .I3(x33_y11)
);

(* keep, dont_touch *)
(* LOC = "X36/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111110000011)
) lut_36_13 (
    .O(x36_y13),
    .I0(x33_y12),
    .I1(1'b0),
    .I2(x34_y8),
    .I3(x34_y18)
);

(* keep, dont_touch *)
(* LOC = "X37/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101000111101)
) lut_37_13 (
    .O(x37_y13),
    .I0(x35_y9),
    .I1(x34_y11),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X38/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011001111001)
) lut_38_13 (
    .O(x38_y13),
    .I0(1'b0),
    .I1(x35_y18),
    .I2(x35_y14),
    .I3(x35_y13)
);

(* keep, dont_touch *)
(* LOC = "X39/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010100100001)
) lut_39_13 (
    .O(x39_y13),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x37_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X40/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110000011010)
) lut_40_13 (
    .O(x40_y13),
    .I0(x38_y18),
    .I1(x38_y13),
    .I2(1'b0),
    .I3(x37_y10)
);

(* keep, dont_touch *)
(* LOC = "X41/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010100100010)
) lut_41_13 (
    .O(x41_y13),
    .I0(x38_y18),
    .I1(1'b0),
    .I2(x39_y18),
    .I3(x38_y13)
);

(* keep, dont_touch *)
(* LOC = "X42/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011100111111)
) lut_42_13 (
    .O(x42_y13),
    .I0(x39_y10),
    .I1(x40_y9),
    .I2(1'b0),
    .I3(x39_y15)
);

(* keep, dont_touch *)
(* LOC = "X43/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010100001011)
) lut_43_13 (
    .O(x43_y13),
    .I0(x40_y15),
    .I1(x40_y18),
    .I2(x41_y11),
    .I3(x40_y13)
);

(* keep, dont_touch *)
(* LOC = "X44/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100010001111)
) lut_44_13 (
    .O(x44_y13),
    .I0(1'b0),
    .I1(x41_y15),
    .I2(x41_y13),
    .I3(x42_y8)
);

(* keep, dont_touch *)
(* LOC = "X45/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110000111101)
) lut_45_13 (
    .O(x45_y13),
    .I0(x43_y16),
    .I1(x42_y9),
    .I2(x43_y12),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X46/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100001001110)
) lut_46_13 (
    .O(x46_y13),
    .I0(x44_y13),
    .I1(x44_y17),
    .I2(x44_y13),
    .I3(x43_y15)
);

(* keep, dont_touch *)
(* LOC = "X47/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000000010110)
) lut_47_13 (
    .O(x47_y13),
    .I0(x44_y13),
    .I1(x45_y18),
    .I2(x44_y11),
    .I3(x45_y13)
);

(* keep, dont_touch *)
(* LOC = "X48/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111010010011)
) lut_48_13 (
    .O(x48_y13),
    .I0(x46_y18),
    .I1(x46_y17),
    .I2(x45_y16),
    .I3(x45_y13)
);

(* keep, dont_touch *)
(* LOC = "X49/Y13" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111000010110)
) lut_49_13 (
    .O(x49_y13),
    .I0(x47_y14),
    .I1(x46_y16),
    .I2(x47_y10),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X0/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010001111011)
) lut_0_14 (
    .O(x0_y14),
    .I0(in4),
    .I1(in9),
    .I2(1'b0),
    .I3(in1)
);

(* keep, dont_touch *)
(* LOC = "X1/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100111010100)
) lut_1_14 (
    .O(x1_y14),
    .I0(in5),
    .I1(in0),
    .I2(1'b0),
    .I3(in7)
);

(* keep, dont_touch *)
(* LOC = "X2/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101000101101)
) lut_2_14 (
    .O(x2_y14),
    .I0(in9),
    .I1(in0),
    .I2(in7),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X3/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100100010100)
) lut_3_14 (
    .O(x3_y14),
    .I0(in8),
    .I1(in8),
    .I2(x1_y14),
    .I3(x1_y13)
);

(* keep, dont_touch *)
(* LOC = "X4/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000100000110)
) lut_4_14 (
    .O(x4_y14),
    .I0(x1_y14),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X5/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100001101100)
) lut_5_14 (
    .O(x5_y14),
    .I0(x2_y9),
    .I1(x3_y18),
    .I2(x2_y14),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X6/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100010010000)
) lut_6_14 (
    .O(x6_y14),
    .I0(x3_y9),
    .I1(x3_y11),
    .I2(x4_y10),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X7/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001011100101)
) lut_7_14 (
    .O(x7_y14),
    .I0(x4_y11),
    .I1(x4_y15),
    .I2(x5_y17),
    .I3(x4_y18)
);

(* keep, dont_touch *)
(* LOC = "X8/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101000101010)
) lut_8_14 (
    .O(x8_y14),
    .I0(x6_y9),
    .I1(x6_y18),
    .I2(x5_y12),
    .I3(x6_y17)
);

(* keep, dont_touch *)
(* LOC = "X9/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100100000000)
) lut_9_14 (
    .O(x9_y14),
    .I0(x6_y9),
    .I1(1'b0),
    .I2(x5_y12),
    .I3(x6_y17)
);

(* keep, dont_touch *)
(* LOC = "X10/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011010101101)
) lut_10_14 (
    .O(x10_y14),
    .I0(x7_y15),
    .I1(x8_y10),
    .I2(1'b0),
    .I3(x8_y18)
);

(* keep, dont_touch *)
(* LOC = "X11/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101010101011)
) lut_11_14 (
    .O(x11_y14),
    .I0(x9_y9),
    .I1(x9_y15),
    .I2(x9_y18),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X12/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010110011010)
) lut_12_14 (
    .O(x12_y14),
    .I0(x9_y15),
    .I1(x10_y11),
    .I2(x9_y17),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X13/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101101101010)
) lut_13_14 (
    .O(x13_y14),
    .I0(x11_y17),
    .I1(x10_y10),
    .I2(1'b0),
    .I3(x10_y19)
);

(* keep, dont_touch *)
(* LOC = "X14/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000011110111)
) lut_14_14 (
    .O(x14_y14),
    .I0(x12_y16),
    .I1(x12_y16),
    .I2(x12_y10),
    .I3(x12_y12)
);

(* keep, dont_touch *)
(* LOC = "X15/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011100110001)
) lut_15_14 (
    .O(x15_y14),
    .I0(x12_y15),
    .I1(x12_y11),
    .I2(x13_y10),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X16/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001001100010)
) lut_16_14 (
    .O(x16_y14),
    .I0(x14_y14),
    .I1(x14_y16),
    .I2(x13_y18),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X17/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111111010011)
) lut_17_14 (
    .O(x17_y14),
    .I0(1'b0),
    .I1(x14_y12),
    .I2(x15_y13),
    .I3(x14_y19)
);

(* keep, dont_touch *)
(* LOC = "X18/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011001110100)
) lut_18_14 (
    .O(x18_y14),
    .I0(x15_y16),
    .I1(1'b0),
    .I2(x15_y12),
    .I3(x15_y10)
);

(* keep, dont_touch *)
(* LOC = "X19/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100111000101)
) lut_19_14 (
    .O(x19_y14),
    .I0(x16_y13),
    .I1(1'b0),
    .I2(x17_y17),
    .I3(x17_y11)
);

(* keep, dont_touch *)
(* LOC = "X20/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111100001111)
) lut_20_14 (
    .O(x20_y14),
    .I0(x18_y15),
    .I1(x17_y17),
    .I2(x18_y14),
    .I3(x18_y19)
);

(* keep, dont_touch *)
(* LOC = "X21/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010101111001)
) lut_21_14 (
    .O(x21_y14),
    .I0(x19_y10),
    .I1(x19_y15),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X22/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001111001110)
) lut_22_14 (
    .O(x22_y14),
    .I0(x19_y16),
    .I1(x20_y14),
    .I2(x20_y19),
    .I3(x19_y19)
);

(* keep, dont_touch *)
(* LOC = "X23/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110111011010)
) lut_23_14 (
    .O(x23_y14),
    .I0(1'b0),
    .I1(x20_y17),
    .I2(x21_y13),
    .I3(x20_y17)
);

(* keep, dont_touch *)
(* LOC = "X24/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101001111110)
) lut_24_14 (
    .O(x24_y14),
    .I0(x22_y16),
    .I1(1'b0),
    .I2(x21_y9),
    .I3(x21_y14)
);

(* keep, dont_touch *)
(* LOC = "X25/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001010101101)
) lut_25_14 (
    .O(x25_y14),
    .I0(1'b0),
    .I1(x23_y18),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X26/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000000111111)
) lut_26_14 (
    .O(x26_y14),
    .I0(x24_y16),
    .I1(1'b0),
    .I2(x23_y10),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X27/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001100010100)
) lut_27_14 (
    .O(x27_y14),
    .I0(x24_y18),
    .I1(x25_y12),
    .I2(x24_y16),
    .I3(x25_y13)
);

(* keep, dont_touch *)
(* LOC = "X28/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111101111100)
) lut_28_14 (
    .O(x28_y14),
    .I0(x25_y15),
    .I1(x26_y13),
    .I2(1'b0),
    .I3(x25_y13)
);

(* keep, dont_touch *)
(* LOC = "X29/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111010101010)
) lut_29_14 (
    .O(x29_y14),
    .I0(x26_y9),
    .I1(1'b0),
    .I2(x26_y12),
    .I3(x27_y11)
);

(* keep, dont_touch *)
(* LOC = "X30/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110011111111)
) lut_30_14 (
    .O(x30_y14),
    .I0(1'b0),
    .I1(x28_y19),
    .I2(x27_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X31/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111101000100)
) lut_31_14 (
    .O(x31_y14),
    .I0(x29_y15),
    .I1(x28_y9),
    .I2(x28_y19),
    .I3(x28_y12)
);

(* keep, dont_touch *)
(* LOC = "X32/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101000110010)
) lut_32_14 (
    .O(x32_y14),
    .I0(x29_y10),
    .I1(x29_y16),
    .I2(x29_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X33/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101000000011)
) lut_33_14 (
    .O(x33_y14),
    .I0(x31_y15),
    .I1(1'b0),
    .I2(x30_y16),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X34/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100000111000)
) lut_34_14 (
    .O(x34_y14),
    .I0(x32_y19),
    .I1(x31_y18),
    .I2(1'b0),
    .I3(x31_y13)
);

(* keep, dont_touch *)
(* LOC = "X35/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010001110000)
) lut_35_14 (
    .O(x35_y14),
    .I0(x32_y10),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x33_y17)
);

(* keep, dont_touch *)
(* LOC = "X36/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000011010000)
) lut_36_14 (
    .O(x36_y14),
    .I0(1'b0),
    .I1(x34_y13),
    .I2(x34_y10),
    .I3(x34_y12)
);

(* keep, dont_touch *)
(* LOC = "X37/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100101000101)
) lut_37_14 (
    .O(x37_y14),
    .I0(x35_y15),
    .I1(x34_y17),
    .I2(x35_y18),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X38/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101111010000)
) lut_38_14 (
    .O(x38_y14),
    .I0(x36_y16),
    .I1(1'b0),
    .I2(x36_y10),
    .I3(x36_y10)
);

(* keep, dont_touch *)
(* LOC = "X39/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100010001001)
) lut_39_14 (
    .O(x39_y14),
    .I0(x37_y18),
    .I1(x37_y13),
    .I2(x37_y16),
    .I3(x37_y19)
);

(* keep, dont_touch *)
(* LOC = "X40/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111111110100)
) lut_40_14 (
    .O(x40_y14),
    .I0(x38_y16),
    .I1(x37_y12),
    .I2(x38_y16),
    .I3(x38_y10)
);

(* keep, dont_touch *)
(* LOC = "X41/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101101010101)
) lut_41_14 (
    .O(x41_y14),
    .I0(1'b0),
    .I1(x39_y9),
    .I2(x38_y12),
    .I3(x38_y10)
);

(* keep, dont_touch *)
(* LOC = "X42/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010101100101)
) lut_42_14 (
    .O(x42_y14),
    .I0(x39_y13),
    .I1(1'b0),
    .I2(x39_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X43/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000000100000)
) lut_43_14 (
    .O(x43_y14),
    .I0(x40_y15),
    .I1(x40_y16),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X44/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001011111011)
) lut_44_14 (
    .O(x44_y14),
    .I0(x41_y16),
    .I1(x42_y12),
    .I2(x41_y18),
    .I3(x42_y16)
);

(* keep, dont_touch *)
(* LOC = "X45/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001010111000)
) lut_45_14 (
    .O(x45_y14),
    .I0(1'b0),
    .I1(x43_y9),
    .I2(x43_y15),
    .I3(x43_y18)
);

(* keep, dont_touch *)
(* LOC = "X46/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100101101110)
) lut_46_14 (
    .O(x46_y14),
    .I0(x43_y19),
    .I1(x43_y16),
    .I2(1'b0),
    .I3(x43_y11)
);

(* keep, dont_touch *)
(* LOC = "X47/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110010000011)
) lut_47_14 (
    .O(x47_y14),
    .I0(1'b0),
    .I1(x45_y14),
    .I2(x44_y11),
    .I3(x44_y17)
);

(* keep, dont_touch *)
(* LOC = "X48/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110001011111)
) lut_48_14 (
    .O(x48_y14),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x45_y12),
    .I3(x46_y10)
);

(* keep, dont_touch *)
(* LOC = "X49/Y14" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010111010111)
) lut_49_14 (
    .O(x49_y14),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x46_y17),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X0/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101101011111)
) lut_0_15 (
    .O(x0_y15),
    .I0(in0),
    .I1(in2),
    .I2(in3),
    .I3(in3)
);

(* keep, dont_touch *)
(* LOC = "X1/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000100001100)
) lut_1_15 (
    .O(x1_y15),
    .I0(in0),
    .I1(in0),
    .I2(in6),
    .I3(in0)
);

(* keep, dont_touch *)
(* LOC = "X2/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011101110111)
) lut_2_15 (
    .O(x2_y15),
    .I0(1'b0),
    .I1(in0),
    .I2(in5),
    .I3(in1)
);

(* keep, dont_touch *)
(* LOC = "X3/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101111100111)
) lut_3_15 (
    .O(x3_y15),
    .I0(1'b0),
    .I1(1'b0),
    .I2(in4),
    .I3(x1_y16)
);

(* keep, dont_touch *)
(* LOC = "X4/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111000011110)
) lut_4_15 (
    .O(x4_y15),
    .I0(x2_y10),
    .I1(x2_y10),
    .I2(x2_y10),
    .I3(x1_y20)
);

(* keep, dont_touch *)
(* LOC = "X5/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000010001011)
) lut_5_15 (
    .O(x5_y15),
    .I0(x3_y14),
    .I1(x3_y10),
    .I2(x3_y16),
    .I3(x2_y17)
);

(* keep, dont_touch *)
(* LOC = "X6/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011001101010)
) lut_6_15 (
    .O(x6_y15),
    .I0(1'b0),
    .I1(x3_y12),
    .I2(1'b0),
    .I3(x4_y19)
);

(* keep, dont_touch *)
(* LOC = "X7/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000100110001)
) lut_7_15 (
    .O(x7_y15),
    .I0(x5_y17),
    .I1(x5_y12),
    .I2(1'b0),
    .I3(x4_y19)
);

(* keep, dont_touch *)
(* LOC = "X8/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000111001110)
) lut_8_15 (
    .O(x8_y15),
    .I0(x6_y12),
    .I1(1'b0),
    .I2(x5_y10),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X9/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000001111110)
) lut_9_15 (
    .O(x9_y15),
    .I0(x7_y14),
    .I1(1'b0),
    .I2(x5_y10),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X10/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100110111000)
) lut_10_15 (
    .O(x10_y15),
    .I0(x8_y15),
    .I1(1'b0),
    .I2(x7_y19),
    .I3(x7_y11)
);

(* keep, dont_touch *)
(* LOC = "X11/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000010111010)
) lut_11_15 (
    .O(x11_y15),
    .I0(1'b0),
    .I1(x9_y18),
    .I2(x8_y18),
    .I3(x8_y20)
);

(* keep, dont_touch *)
(* LOC = "X12/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001001101100)
) lut_12_15 (
    .O(x12_y15),
    .I0(x10_y17),
    .I1(1'b0),
    .I2(x9_y15),
    .I3(x9_y17)
);

(* keep, dont_touch *)
(* LOC = "X13/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010011001001)
) lut_13_15 (
    .O(x13_y15),
    .I0(x10_y10),
    .I1(x10_y20),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X14/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100001101011)
) lut_14_15 (
    .O(x14_y15),
    .I0(1'b0),
    .I1(x11_y18),
    .I2(1'b0),
    .I3(x11_y12)
);

(* keep, dont_touch *)
(* LOC = "X15/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101010010101)
) lut_15_15 (
    .O(x15_y15),
    .I0(x12_y10),
    .I1(x13_y16),
    .I2(x13_y18),
    .I3(x12_y12)
);

(* keep, dont_touch *)
(* LOC = "X16/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001101111011)
) lut_16_15 (
    .O(x16_y15),
    .I0(x13_y10),
    .I1(x13_y17),
    .I2(x13_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X17/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111011010100)
) lut_17_15 (
    .O(x17_y15),
    .I0(x14_y10),
    .I1(x14_y14),
    .I2(x14_y19),
    .I3(x15_y18)
);

(* keep, dont_touch *)
(* LOC = "X18/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011000101001)
) lut_18_15 (
    .O(x18_y15),
    .I0(1'b0),
    .I1(x15_y13),
    .I2(x16_y20),
    .I3(x16_y20)
);

(* keep, dont_touch *)
(* LOC = "X19/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010010011100)
) lut_19_15 (
    .O(x19_y15),
    .I0(x17_y11),
    .I1(x17_y11),
    .I2(x16_y14),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X20/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010111100110)
) lut_20_15 (
    .O(x20_y15),
    .I0(x18_y10),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X21/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110011111011)
) lut_21_15 (
    .O(x21_y15),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x19_y19)
);

(* keep, dont_touch *)
(* LOC = "X22/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100010110010)
) lut_22_15 (
    .O(x22_y15),
    .I0(x19_y13),
    .I1(x20_y16),
    .I2(x19_y17),
    .I3(x20_y14)
);

(* keep, dont_touch *)
(* LOC = "X23/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100101001110)
) lut_23_15 (
    .O(x23_y15),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x21_y13),
    .I3(x20_y11)
);

(* keep, dont_touch *)
(* LOC = "X24/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010011000111)
) lut_24_15 (
    .O(x24_y15),
    .I0(1'b0),
    .I1(x21_y16),
    .I2(x21_y15),
    .I3(x21_y16)
);

(* keep, dont_touch *)
(* LOC = "X25/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001010011101)
) lut_25_15 (
    .O(x25_y15),
    .I0(x23_y15),
    .I1(x23_y16),
    .I2(x23_y16),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X26/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101110011110)
) lut_26_15 (
    .O(x26_y15),
    .I0(x23_y20),
    .I1(x23_y13),
    .I2(1'b0),
    .I3(x24_y12)
);

(* keep, dont_touch *)
(* LOC = "X27/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011001110101)
) lut_27_15 (
    .O(x27_y15),
    .I0(x24_y12),
    .I1(x25_y11),
    .I2(x25_y15),
    .I3(x25_y13)
);

(* keep, dont_touch *)
(* LOC = "X28/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011000010001)
) lut_28_15 (
    .O(x28_y15),
    .I0(1'b0),
    .I1(x26_y11),
    .I2(x25_y10),
    .I3(x26_y14)
);

(* keep, dont_touch *)
(* LOC = "X29/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011000001001)
) lut_29_15 (
    .O(x29_y15),
    .I0(x26_y18),
    .I1(x27_y11),
    .I2(x26_y12),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X30/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110111010100)
) lut_30_15 (
    .O(x30_y15),
    .I0(1'b0),
    .I1(x27_y10),
    .I2(1'b0),
    .I3(x28_y10)
);

(* keep, dont_touch *)
(* LOC = "X31/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100101101011)
) lut_31_15 (
    .O(x31_y15),
    .I0(1'b0),
    .I1(x29_y18),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X32/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100101000001)
) lut_32_15 (
    .O(x32_y15),
    .I0(1'b0),
    .I1(x30_y19),
    .I2(x30_y19),
    .I3(x29_y17)
);

(* keep, dont_touch *)
(* LOC = "X33/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100001111110)
) lut_33_15 (
    .O(x33_y15),
    .I0(x31_y19),
    .I1(x30_y10),
    .I2(x31_y16),
    .I3(x30_y10)
);

(* keep, dont_touch *)
(* LOC = "X34/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011000111010)
) lut_34_15 (
    .O(x34_y15),
    .I0(1'b0),
    .I1(x32_y19),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X35/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000100010011)
) lut_35_15 (
    .O(x35_y15),
    .I0(x32_y15),
    .I1(x32_y14),
    .I2(x33_y15),
    .I3(x32_y14)
);

(* keep, dont_touch *)
(* LOC = "X36/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011011100000)
) lut_36_15 (
    .O(x36_y15),
    .I0(x33_y12),
    .I1(x34_y15),
    .I2(1'b0),
    .I3(x34_y14)
);

(* keep, dont_touch *)
(* LOC = "X37/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101000010101)
) lut_37_15 (
    .O(x37_y15),
    .I0(x34_y17),
    .I1(x35_y14),
    .I2(1'b0),
    .I3(x34_y15)
);

(* keep, dont_touch *)
(* LOC = "X38/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110001000000)
) lut_38_15 (
    .O(x38_y15),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x35_y12)
);

(* keep, dont_touch *)
(* LOC = "X39/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000100110001)
) lut_39_15 (
    .O(x39_y15),
    .I0(x37_y15),
    .I1(x37_y20),
    .I2(1'b0),
    .I3(x36_y19)
);

(* keep, dont_touch *)
(* LOC = "X40/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001100011000)
) lut_40_15 (
    .O(x40_y15),
    .I0(x37_y13),
    .I1(x38_y18),
    .I2(x38_y19),
    .I3(x37_y19)
);

(* keep, dont_touch *)
(* LOC = "X41/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111000110111)
) lut_41_15 (
    .O(x41_y15),
    .I0(1'b0),
    .I1(x39_y19),
    .I2(x38_y16),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X42/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000101001101)
) lut_42_15 (
    .O(x42_y15),
    .I0(x39_y19),
    .I1(x40_y15),
    .I2(x40_y15),
    .I3(x40_y14)
);

(* keep, dont_touch *)
(* LOC = "X43/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011100010001)
) lut_43_15 (
    .O(x43_y15),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x40_y14),
    .I3(x40_y10)
);

(* keep, dont_touch *)
(* LOC = "X44/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000011001111)
) lut_44_15 (
    .O(x44_y15),
    .I0(x41_y20),
    .I1(x41_y12),
    .I2(1'b0),
    .I3(x42_y20)
);

(* keep, dont_touch *)
(* LOC = "X45/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001101000111)
) lut_45_15 (
    .O(x45_y15),
    .I0(x43_y11),
    .I1(x42_y15),
    .I2(x42_y20),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X46/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111011000101)
) lut_46_15 (
    .O(x46_y15),
    .I0(1'b0),
    .I1(x43_y19),
    .I2(x43_y18),
    .I3(x43_y19)
);

(* keep, dont_touch *)
(* LOC = "X47/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110100111110)
) lut_47_15 (
    .O(x47_y15),
    .I0(x44_y16),
    .I1(x45_y12),
    .I2(x44_y20),
    .I3(x44_y15)
);

(* keep, dont_touch *)
(* LOC = "X48/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101001111110)
) lut_48_15 (
    .O(x48_y15),
    .I0(x45_y18),
    .I1(x45_y17),
    .I2(x45_y19),
    .I3(x45_y13)
);

(* keep, dont_touch *)
(* LOC = "X49/Y15" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000101011000)
) lut_49_15 (
    .O(x49_y15),
    .I0(x47_y16),
    .I1(x47_y16),
    .I2(x46_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X0/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001010001011)
) lut_0_16 (
    .O(x0_y16),
    .I0(in1),
    .I1(in2),
    .I2(in6),
    .I3(in6)
);

(* keep, dont_touch *)
(* LOC = "X1/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011001010011)
) lut_1_16 (
    .O(x1_y16),
    .I0(in2),
    .I1(in4),
    .I2(in1),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X2/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110010000101)
) lut_2_16 (
    .O(x2_y16),
    .I0(in1),
    .I1(1'b0),
    .I2(in2),
    .I3(in1)
);

(* keep, dont_touch *)
(* LOC = "X3/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111000111111)
) lut_3_16 (
    .O(x3_y16),
    .I0(1'b0),
    .I1(1'b0),
    .I2(in0),
    .I3(in1)
);

(* keep, dont_touch *)
(* LOC = "X4/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010101111110)
) lut_4_16 (
    .O(x4_y16),
    .I0(1'b0),
    .I1(x1_y20),
    .I2(1'b0),
    .I3(x2_y20)
);

(* keep, dont_touch *)
(* LOC = "X5/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100010100111)
) lut_5_16 (
    .O(x5_y16),
    .I0(x2_y19),
    .I1(x2_y19),
    .I2(1'b0),
    .I3(x2_y11)
);

(* keep, dont_touch *)
(* LOC = "X6/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011111000111)
) lut_6_16 (
    .O(x6_y16),
    .I0(x3_y20),
    .I1(x4_y17),
    .I2(x4_y17),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X7/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110100011111)
) lut_7_16 (
    .O(x7_y16),
    .I0(x4_y13),
    .I1(x5_y20),
    .I2(1'b0),
    .I3(x5_y17)
);

(* keep, dont_touch *)
(* LOC = "X8/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010100010100)
) lut_8_16 (
    .O(x8_y16),
    .I0(x6_y19),
    .I1(x6_y15),
    .I2(x5_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X9/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001110000011)
) lut_9_16 (
    .O(x9_y16),
    .I0(x6_y16),
    .I1(1'b0),
    .I2(x5_y11),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X10/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000000110111)
) lut_10_16 (
    .O(x10_y16),
    .I0(x7_y13),
    .I1(x8_y15),
    .I2(x8_y15),
    .I3(x7_y11)
);

(* keep, dont_touch *)
(* LOC = "X11/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100001100001)
) lut_11_16 (
    .O(x11_y16),
    .I0(x8_y20),
    .I1(x8_y20),
    .I2(x8_y15),
    .I3(x8_y18)
);

(* keep, dont_touch *)
(* LOC = "X12/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100110100000)
) lut_12_16 (
    .O(x12_y16),
    .I0(x10_y14),
    .I1(x9_y13),
    .I2(x9_y15),
    .I3(x10_y19)
);

(* keep, dont_touch *)
(* LOC = "X13/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010100001100)
) lut_13_16 (
    .O(x13_y16),
    .I0(1'b0),
    .I1(x11_y11),
    .I2(x10_y20),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X14/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111101011000)
) lut_14_16 (
    .O(x14_y16),
    .I0(1'b0),
    .I1(x12_y16),
    .I2(x11_y16),
    .I3(x11_y21)
);

(* keep, dont_touch *)
(* LOC = "X15/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000001010000)
) lut_15_16 (
    .O(x15_y16),
    .I0(1'b0),
    .I1(x12_y16),
    .I2(1'b0),
    .I3(x13_y14)
);

(* keep, dont_touch *)
(* LOC = "X16/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001000110000)
) lut_16_16 (
    .O(x16_y16),
    .I0(x13_y19),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X17/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101001111100)
) lut_17_16 (
    .O(x17_y16),
    .I0(x14_y18),
    .I1(x15_y21),
    .I2(x15_y20),
    .I3(x15_y19)
);

(* keep, dont_touch *)
(* LOC = "X18/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001000001000)
) lut_18_16 (
    .O(x18_y16),
    .I0(x16_y18),
    .I1(x15_y14),
    .I2(x15_y17),
    .I3(x16_y18)
);

(* keep, dont_touch *)
(* LOC = "X19/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000101000011)
) lut_19_16 (
    .O(x19_y16),
    .I0(x17_y11),
    .I1(x16_y19),
    .I2(1'b0),
    .I3(x17_y14)
);

(* keep, dont_touch *)
(* LOC = "X20/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100010010001)
) lut_20_16 (
    .O(x20_y16),
    .I0(x17_y18),
    .I1(x17_y21),
    .I2(x18_y14),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X21/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001101011011)
) lut_21_16 (
    .O(x21_y16),
    .I0(x18_y12),
    .I1(x19_y11),
    .I2(x19_y19),
    .I3(x18_y11)
);

(* keep, dont_touch *)
(* LOC = "X22/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011001101010)
) lut_22_16 (
    .O(x22_y16),
    .I0(x20_y17),
    .I1(x19_y16),
    .I2(x19_y20),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X23/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011000001000)
) lut_23_16 (
    .O(x23_y16),
    .I0(x21_y19),
    .I1(x21_y19),
    .I2(x21_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X24/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011101011110)
) lut_24_16 (
    .O(x24_y16),
    .I0(1'b0),
    .I1(x22_y17),
    .I2(1'b0),
    .I3(x22_y14)
);

(* keep, dont_touch *)
(* LOC = "X25/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011101011001)
) lut_25_16 (
    .O(x25_y16),
    .I0(x23_y19),
    .I1(x23_y19),
    .I2(x22_y11),
    .I3(x22_y16)
);

(* keep, dont_touch *)
(* LOC = "X26/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110101111110)
) lut_26_16 (
    .O(x26_y16),
    .I0(x23_y21),
    .I1(x23_y13),
    .I2(x24_y17),
    .I3(x23_y11)
);

(* keep, dont_touch *)
(* LOC = "X27/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000000000001)
) lut_27_16 (
    .O(x27_y16),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x25_y21),
    .I3(x24_y14)
);

(* keep, dont_touch *)
(* LOC = "X28/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100101001000)
) lut_28_16 (
    .O(x28_y16),
    .I0(x26_y16),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x25_y11)
);

(* keep, dont_touch *)
(* LOC = "X29/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100110010111)
) lut_29_16 (
    .O(x29_y16),
    .I0(1'b0),
    .I1(x27_y20),
    .I2(x26_y12),
    .I3(x26_y16)
);

(* keep, dont_touch *)
(* LOC = "X30/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010101000011)
) lut_30_16 (
    .O(x30_y16),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x28_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X31/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000110011011)
) lut_31_16 (
    .O(x31_y16),
    .I0(x29_y12),
    .I1(1'b0),
    .I2(x28_y11),
    .I3(x29_y11)
);

(* keep, dont_touch *)
(* LOC = "X32/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111100011011)
) lut_32_16 (
    .O(x32_y16),
    .I0(x30_y18),
    .I1(1'b0),
    .I2(x30_y11),
    .I3(x30_y13)
);

(* keep, dont_touch *)
(* LOC = "X33/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000001110010)
) lut_33_16 (
    .O(x33_y16),
    .I0(x30_y19),
    .I1(1'b0),
    .I2(x31_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X34/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100111000101)
) lut_34_16 (
    .O(x34_y16),
    .I0(x31_y14),
    .I1(x32_y16),
    .I2(x31_y15),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X35/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011111001000)
) lut_35_16 (
    .O(x35_y16),
    .I0(x33_y18),
    .I1(x32_y11),
    .I2(x32_y17),
    .I3(x33_y20)
);

(* keep, dont_touch *)
(* LOC = "X36/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111010111111)
) lut_36_16 (
    .O(x36_y16),
    .I0(1'b0),
    .I1(x34_y16),
    .I2(x34_y12),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X37/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010110101101)
) lut_37_16 (
    .O(x37_y16),
    .I0(x35_y16),
    .I1(x35_y19),
    .I2(1'b0),
    .I3(x34_y16)
);

(* keep, dont_touch *)
(* LOC = "X38/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001011000000)
) lut_38_16 (
    .O(x38_y16),
    .I0(x36_y21),
    .I1(x36_y16),
    .I2(x36_y19),
    .I3(x35_y12)
);

(* keep, dont_touch *)
(* LOC = "X39/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000110110011)
) lut_39_16 (
    .O(x39_y16),
    .I0(1'b0),
    .I1(x37_y16),
    .I2(1'b0),
    .I3(x37_y12)
);

(* keep, dont_touch *)
(* LOC = "X40/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110010000100)
) lut_40_16 (
    .O(x40_y16),
    .I0(x38_y11),
    .I1(x37_y18),
    .I2(1'b0),
    .I3(x38_y20)
);

(* keep, dont_touch *)
(* LOC = "X41/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001111101000)
) lut_41_16 (
    .O(x41_y16),
    .I0(x39_y14),
    .I1(x39_y15),
    .I2(x39_y11),
    .I3(x39_y16)
);

(* keep, dont_touch *)
(* LOC = "X42/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001101111100)
) lut_42_16 (
    .O(x42_y16),
    .I0(x40_y16),
    .I1(x39_y15),
    .I2(x40_y15),
    .I3(x40_y18)
);

(* keep, dont_touch *)
(* LOC = "X43/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001110110001)
) lut_43_16 (
    .O(x43_y16),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x41_y11),
    .I3(x40_y12)
);

(* keep, dont_touch *)
(* LOC = "X44/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101100000100)
) lut_44_16 (
    .O(x44_y16),
    .I0(x41_y17),
    .I1(1'b0),
    .I2(x42_y19),
    .I3(x42_y21)
);

(* keep, dont_touch *)
(* LOC = "X45/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110111111010)
) lut_45_16 (
    .O(x45_y16),
    .I0(x42_y13),
    .I1(1'b0),
    .I2(x42_y18),
    .I3(x42_y15)
);

(* keep, dont_touch *)
(* LOC = "X46/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011010100010)
) lut_46_16 (
    .O(x46_y16),
    .I0(x43_y13),
    .I1(x43_y20),
    .I2(x44_y19),
    .I3(x43_y16)
);

(* keep, dont_touch *)
(* LOC = "X47/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100101101011)
) lut_47_16 (
    .O(x47_y16),
    .I0(x45_y12),
    .I1(x44_y11),
    .I2(1'b0),
    .I3(x44_y15)
);

(* keep, dont_touch *)
(* LOC = "X48/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011111000010)
) lut_48_16 (
    .O(x48_y16),
    .I0(x46_y13),
    .I1(x45_y19),
    .I2(x46_y12),
    .I3(x46_y15)
);

(* keep, dont_touch *)
(* LOC = "X49/Y16" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100101010101)
) lut_49_16 (
    .O(x49_y16),
    .I0(x46_y12),
    .I1(x47_y20),
    .I2(x47_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X0/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111000011011)
) lut_0_17 (
    .O(x0_y17),
    .I0(1'b0),
    .I1(1'b0),
    .I2(in7),
    .I3(in4)
);

(* keep, dont_touch *)
(* LOC = "X1/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111111111010)
) lut_1_17 (
    .O(x1_y17),
    .I0(in0),
    .I1(in0),
    .I2(in7),
    .I3(in2)
);

(* keep, dont_touch *)
(* LOC = "X2/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000110101110)
) lut_2_17 (
    .O(x2_y17),
    .I0(1'b0),
    .I1(in6),
    .I2(in2),
    .I3(in7)
);

(* keep, dont_touch *)
(* LOC = "X3/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011101001111)
) lut_3_17 (
    .O(x3_y17),
    .I0(x1_y12),
    .I1(in0),
    .I2(in7),
    .I3(x1_y18)
);

(* keep, dont_touch *)
(* LOC = "X4/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110101111110)
) lut_4_17 (
    .O(x4_y17),
    .I0(1'b0),
    .I1(x2_y17),
    .I2(1'b0),
    .I3(x1_y17)
);

(* keep, dont_touch *)
(* LOC = "X5/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000001110011)
) lut_5_17 (
    .O(x5_y17),
    .I0(x3_y19),
    .I1(x2_y14),
    .I2(x3_y17),
    .I3(x3_y15)
);

(* keep, dont_touch *)
(* LOC = "X6/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010100111010)
) lut_6_17 (
    .O(x6_y17),
    .I0(x3_y12),
    .I1(1'b0),
    .I2(x4_y21),
    .I3(x3_y15)
);

(* keep, dont_touch *)
(* LOC = "X7/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100100011110)
) lut_7_17 (
    .O(x7_y17),
    .I0(x5_y15),
    .I1(x5_y18),
    .I2(x5_y21),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X8/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100001001110)
) lut_8_17 (
    .O(x8_y17),
    .I0(x5_y20),
    .I1(x5_y18),
    .I2(x6_y13),
    .I3(x5_y20)
);

(* keep, dont_touch *)
(* LOC = "X9/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111011000001)
) lut_9_17 (
    .O(x9_y17),
    .I0(x6_y14),
    .I1(x6_y14),
    .I2(x6_y13),
    .I3(x5_y20)
);

(* keep, dont_touch *)
(* LOC = "X10/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000001000010)
) lut_10_17 (
    .O(x10_y17),
    .I0(x7_y15),
    .I1(1'b0),
    .I2(x8_y22),
    .I3(x8_y19)
);

(* keep, dont_touch *)
(* LOC = "X11/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000111000010)
) lut_11_17 (
    .O(x11_y17),
    .I0(1'b0),
    .I1(x9_y15),
    .I2(x8_y13),
    .I3(x9_y12)
);

(* keep, dont_touch *)
(* LOC = "X12/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010001110111)
) lut_12_17 (
    .O(x12_y17),
    .I0(1'b0),
    .I1(x10_y14),
    .I2(x9_y22),
    .I3(x10_y20)
);

(* keep, dont_touch *)
(* LOC = "X13/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011011001000)
) lut_13_17 (
    .O(x13_y17),
    .I0(x11_y15),
    .I1(x10_y14),
    .I2(x10_y19),
    .I3(x11_y12)
);

(* keep, dont_touch *)
(* LOC = "X14/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011010000100)
) lut_14_17 (
    .O(x14_y17),
    .I0(1'b0),
    .I1(x12_y22),
    .I2(x11_y14),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X15/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101111000001)
) lut_15_17 (
    .O(x15_y17),
    .I0(x12_y18),
    .I1(1'b0),
    .I2(x13_y21),
    .I3(x12_y21)
);

(* keep, dont_touch *)
(* LOC = "X16/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011101111111)
) lut_16_17 (
    .O(x16_y17),
    .I0(x13_y15),
    .I1(x14_y13),
    .I2(x14_y21),
    .I3(x14_y21)
);

(* keep, dont_touch *)
(* LOC = "X17/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011000111000)
) lut_17_17 (
    .O(x17_y17),
    .I0(x14_y14),
    .I1(x15_y19),
    .I2(x15_y16),
    .I3(x15_y21)
);

(* keep, dont_touch *)
(* LOC = "X18/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100100101001)
) lut_18_17 (
    .O(x18_y17),
    .I0(x15_y22),
    .I1(1'b0),
    .I2(x16_y21),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X19/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110000001010)
) lut_19_17 (
    .O(x19_y17),
    .I0(1'b0),
    .I1(x16_y15),
    .I2(x16_y17),
    .I3(x17_y16)
);

(* keep, dont_touch *)
(* LOC = "X20/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110110010100)
) lut_20_17 (
    .O(x20_y17),
    .I0(1'b0),
    .I1(x18_y15),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X21/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011111110001)
) lut_21_17 (
    .O(x21_y17),
    .I0(x18_y13),
    .I1(x19_y22),
    .I2(x18_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X22/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011101010011)
) lut_22_17 (
    .O(x22_y17),
    .I0(x19_y18),
    .I1(x19_y13),
    .I2(x20_y16),
    .I3(x20_y22)
);

(* keep, dont_touch *)
(* LOC = "X23/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111100001000)
) lut_23_17 (
    .O(x23_y17),
    .I0(x20_y12),
    .I1(x21_y16),
    .I2(x21_y14),
    .I3(x20_y15)
);

(* keep, dont_touch *)
(* LOC = "X24/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001000101011)
) lut_24_17 (
    .O(x24_y17),
    .I0(1'b0),
    .I1(x22_y19),
    .I2(1'b0),
    .I3(x22_y22)
);

(* keep, dont_touch *)
(* LOC = "X25/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000001110011)
) lut_25_17 (
    .O(x25_y17),
    .I0(1'b0),
    .I1(x22_y12),
    .I2(1'b0),
    .I3(x22_y14)
);

(* keep, dont_touch *)
(* LOC = "X26/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001000011101)
) lut_26_17 (
    .O(x26_y17),
    .I0(x24_y13),
    .I1(x24_y16),
    .I2(x23_y17),
    .I3(x24_y19)
);

(* keep, dont_touch *)
(* LOC = "X27/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010011011001)
) lut_27_17 (
    .O(x27_y17),
    .I0(x25_y16),
    .I1(x25_y19),
    .I2(x25_y13),
    .I3(x25_y16)
);

(* keep, dont_touch *)
(* LOC = "X28/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000100000100)
) lut_28_17 (
    .O(x28_y17),
    .I0(x26_y22),
    .I1(x26_y20),
    .I2(1'b0),
    .I3(x26_y18)
);

(* keep, dont_touch *)
(* LOC = "X29/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001010100000)
) lut_29_17 (
    .O(x29_y17),
    .I0(x27_y22),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X30/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101101001101)
) lut_30_17 (
    .O(x30_y17),
    .I0(x28_y13),
    .I1(x28_y15),
    .I2(1'b0),
    .I3(x28_y21)
);

(* keep, dont_touch *)
(* LOC = "X31/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101001001001)
) lut_31_17 (
    .O(x31_y17),
    .I0(x29_y16),
    .I1(1'b0),
    .I2(x28_y19),
    .I3(x29_y13)
);

(* keep, dont_touch *)
(* LOC = "X32/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110101101011)
) lut_32_17 (
    .O(x32_y17),
    .I0(x29_y22),
    .I1(x30_y14),
    .I2(1'b0),
    .I3(x30_y21)
);

(* keep, dont_touch *)
(* LOC = "X33/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101011011111)
) lut_33_17 (
    .O(x33_y17),
    .I0(x31_y14),
    .I1(x31_y22),
    .I2(x31_y18),
    .I3(x30_y14)
);

(* keep, dont_touch *)
(* LOC = "X34/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010010010111)
) lut_34_17 (
    .O(x34_y17),
    .I0(x31_y16),
    .I1(x32_y16),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X35/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011111001101)
) lut_35_17 (
    .O(x35_y17),
    .I0(x33_y14),
    .I1(x32_y16),
    .I2(x33_y20),
    .I3(x33_y21)
);

(* keep, dont_touch *)
(* LOC = "X36/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111100000101)
) lut_36_17 (
    .O(x36_y17),
    .I0(x34_y17),
    .I1(x33_y16),
    .I2(x33_y18),
    .I3(x33_y20)
);

(* keep, dont_touch *)
(* LOC = "X37/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101011010011)
) lut_37_17 (
    .O(x37_y17),
    .I0(x35_y16),
    .I1(x35_y17),
    .I2(x34_y18),
    .I3(x35_y18)
);

(* keep, dont_touch *)
(* LOC = "X38/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001101011111)
) lut_38_17 (
    .O(x38_y17),
    .I0(x36_y21),
    .I1(1'b0),
    .I2(x35_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X39/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011010111111)
) lut_39_17 (
    .O(x39_y17),
    .I0(x37_y14),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x36_y16)
);

(* keep, dont_touch *)
(* LOC = "X40/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101001100010)
) lut_40_17 (
    .O(x40_y17),
    .I0(x38_y16),
    .I1(x37_y13),
    .I2(x38_y21),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X41/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010011010000)
) lut_41_17 (
    .O(x41_y17),
    .I0(x38_y13),
    .I1(x39_y18),
    .I2(x38_y17),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X42/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000001011010)
) lut_42_17 (
    .O(x42_y17),
    .I0(1'b0),
    .I1(x39_y22),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X43/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000110001101)
) lut_43_17 (
    .O(x43_y17),
    .I0(x40_y15),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X44/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011111001110)
) lut_44_17 (
    .O(x44_y17),
    .I0(1'b0),
    .I1(x42_y12),
    .I2(x42_y15),
    .I3(x41_y18)
);

(* keep, dont_touch *)
(* LOC = "X45/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110101001100)
) lut_45_17 (
    .O(x45_y17),
    .I0(x42_y18),
    .I1(x42_y15),
    .I2(x43_y21),
    .I3(x42_y16)
);

(* keep, dont_touch *)
(* LOC = "X46/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010111101000)
) lut_46_17 (
    .O(x46_y17),
    .I0(1'b0),
    .I1(x44_y20),
    .I2(x44_y12),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X47/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011011010100)
) lut_47_17 (
    .O(x47_y17),
    .I0(x44_y12),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X48/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101000100010)
) lut_48_17 (
    .O(x48_y17),
    .I0(x46_y18),
    .I1(x45_y21),
    .I2(x45_y16),
    .I3(x45_y17)
);

(* keep, dont_touch *)
(* LOC = "X49/Y17" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101111011011)
) lut_49_17 (
    .O(x49_y17),
    .I0(x47_y17),
    .I1(1'b0),
    .I2(x47_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X0/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111010001101)
) lut_0_18 (
    .O(x0_y18),
    .I0(1'b0),
    .I1(in4),
    .I2(in3),
    .I3(in9)
);

(* keep, dont_touch *)
(* LOC = "X1/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011001000011)
) lut_1_18 (
    .O(x1_y18),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X2/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001111111010)
) lut_2_18 (
    .O(x2_y18),
    .I0(in5),
    .I1(in3),
    .I2(1'b0),
    .I3(in8)
);

(* keep, dont_touch *)
(* LOC = "X3/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101011110000)
) lut_3_18 (
    .O(x3_y18),
    .I0(in9),
    .I1(in2),
    .I2(x1_y22),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X4/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010001100010)
) lut_4_18 (
    .O(x4_y18),
    .I0(1'b0),
    .I1(x2_y20),
    .I2(x2_y23),
    .I3(x2_y22)
);

(* keep, dont_touch *)
(* LOC = "X5/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000101011010)
) lut_5_18 (
    .O(x5_y18),
    .I0(x3_y22),
    .I1(x2_y18),
    .I2(x3_y20),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X6/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000101110100)
) lut_6_18 (
    .O(x6_y18),
    .I0(x4_y19),
    .I1(x4_y19),
    .I2(x4_y20),
    .I3(x4_y23)
);

(* keep, dont_touch *)
(* LOC = "X7/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001110000000)
) lut_7_18 (
    .O(x7_y18),
    .I0(1'b0),
    .I1(x4_y16),
    .I2(1'b0),
    .I3(x4_y13)
);

(* keep, dont_touch *)
(* LOC = "X8/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011110100001)
) lut_8_18 (
    .O(x8_y18),
    .I0(x6_y18),
    .I1(x5_y17),
    .I2(x6_y15),
    .I3(x6_y22)
);

(* keep, dont_touch *)
(* LOC = "X9/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101100010110)
) lut_9_18 (
    .O(x9_y18),
    .I0(x7_y22),
    .I1(x6_y21),
    .I2(x6_y15),
    .I3(x6_y22)
);

(* keep, dont_touch *)
(* LOC = "X10/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111100111001)
) lut_10_18 (
    .O(x10_y18),
    .I0(x7_y13),
    .I1(1'b0),
    .I2(x8_y23),
    .I3(x7_y13)
);

(* keep, dont_touch *)
(* LOC = "X11/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101010110110)
) lut_11_18 (
    .O(x11_y18),
    .I0(x9_y13),
    .I1(x9_y18),
    .I2(x8_y18),
    .I3(x9_y16)
);

(* keep, dont_touch *)
(* LOC = "X12/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111010010010)
) lut_12_18 (
    .O(x12_y18),
    .I0(x10_y13),
    .I1(x9_y19),
    .I2(x9_y13),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X13/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110000100100)
) lut_13_18 (
    .O(x13_y18),
    .I0(x10_y21),
    .I1(x10_y21),
    .I2(x11_y22),
    .I3(x10_y14)
);

(* keep, dont_touch *)
(* LOC = "X14/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110010100000)
) lut_14_18 (
    .O(x14_y18),
    .I0(x11_y14),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x12_y22)
);

(* keep, dont_touch *)
(* LOC = "X15/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100001000010)
) lut_15_18 (
    .O(x15_y18),
    .I0(1'b0),
    .I1(x12_y20),
    .I2(x12_y22),
    .I3(x12_y15)
);

(* keep, dont_touch *)
(* LOC = "X16/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000110110011)
) lut_16_18 (
    .O(x16_y18),
    .I0(x13_y20),
    .I1(1'b0),
    .I2(x13_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X17/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001000011110)
) lut_17_18 (
    .O(x17_y18),
    .I0(x14_y15),
    .I1(x15_y14),
    .I2(x14_y14),
    .I3(x14_y16)
);

(* keep, dont_touch *)
(* LOC = "X18/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101011110010)
) lut_18_18 (
    .O(x18_y18),
    .I0(1'b0),
    .I1(x15_y17),
    .I2(x15_y16),
    .I3(x16_y14)
);

(* keep, dont_touch *)
(* LOC = "X19/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111011000110)
) lut_19_18 (
    .O(x19_y18),
    .I0(x17_y21),
    .I1(x17_y20),
    .I2(1'b0),
    .I3(x16_y23)
);

(* keep, dont_touch *)
(* LOC = "X20/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011100100101)
) lut_20_18 (
    .O(x20_y18),
    .I0(x18_y13),
    .I1(x17_y23),
    .I2(x18_y17),
    .I3(x17_y22)
);

(* keep, dont_touch *)
(* LOC = "X21/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011111001110)
) lut_21_18 (
    .O(x21_y18),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x18_y22)
);

(* keep, dont_touch *)
(* LOC = "X22/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111111010101)
) lut_22_18 (
    .O(x22_y18),
    .I0(x19_y23),
    .I1(1'b0),
    .I2(x19_y15),
    .I3(x19_y14)
);

(* keep, dont_touch *)
(* LOC = "X23/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111011101010)
) lut_23_18 (
    .O(x23_y18),
    .I0(x21_y16),
    .I1(x21_y15),
    .I2(x21_y22),
    .I3(x21_y19)
);

(* keep, dont_touch *)
(* LOC = "X24/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110001100100)
) lut_24_18 (
    .O(x24_y18),
    .I0(x22_y14),
    .I1(x22_y17),
    .I2(x21_y21),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X25/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110110000001)
) lut_25_18 (
    .O(x25_y18),
    .I0(x22_y21),
    .I1(1'b0),
    .I2(x23_y20),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X26/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010000100111)
) lut_26_18 (
    .O(x26_y18),
    .I0(x24_y15),
    .I1(x24_y17),
    .I2(x23_y23),
    .I3(x24_y18)
);

(* keep, dont_touch *)
(* LOC = "X27/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011101010001)
) lut_27_18 (
    .O(x27_y18),
    .I0(x25_y20),
    .I1(x25_y23),
    .I2(x24_y16),
    .I3(x24_y17)
);

(* keep, dont_touch *)
(* LOC = "X28/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111101001110)
) lut_28_18 (
    .O(x28_y18),
    .I0(1'b0),
    .I1(x25_y21),
    .I2(x26_y13),
    .I3(x26_y14)
);

(* keep, dont_touch *)
(* LOC = "X29/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001110010000)
) lut_29_18 (
    .O(x29_y18),
    .I0(1'b0),
    .I1(x26_y16),
    .I2(x27_y21),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X30/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101011111100)
) lut_30_18 (
    .O(x30_y18),
    .I0(x27_y16),
    .I1(x28_y21),
    .I2(x27_y23),
    .I3(x27_y13)
);

(* keep, dont_touch *)
(* LOC = "X31/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001011010111)
) lut_31_18 (
    .O(x31_y18),
    .I0(x28_y15),
    .I1(1'b0),
    .I2(x29_y23),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X32/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100010101011)
) lut_32_18 (
    .O(x32_y18),
    .I0(x29_y18),
    .I1(x29_y17),
    .I2(x30_y23),
    .I3(x29_y21)
);

(* keep, dont_touch *)
(* LOC = "X33/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101010000011)
) lut_33_18 (
    .O(x33_y18),
    .I0(x31_y19),
    .I1(1'b0),
    .I2(x30_y18),
    .I3(x30_y14)
);

(* keep, dont_touch *)
(* LOC = "X34/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111000110100)
) lut_34_18 (
    .O(x34_y18),
    .I0(x32_y18),
    .I1(x31_y21),
    .I2(x32_y19),
    .I3(x31_y18)
);

(* keep, dont_touch *)
(* LOC = "X35/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110110000000)
) lut_35_18 (
    .O(x35_y18),
    .I0(1'b0),
    .I1(x32_y17),
    .I2(x33_y13),
    .I3(x33_y18)
);

(* keep, dont_touch *)
(* LOC = "X36/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110101110000)
) lut_36_18 (
    .O(x36_y18),
    .I0(x33_y21),
    .I1(x33_y16),
    .I2(x33_y15),
    .I3(x34_y18)
);

(* keep, dont_touch *)
(* LOC = "X37/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010010101101)
) lut_37_18 (
    .O(x37_y18),
    .I0(x35_y18),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X38/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100100110101)
) lut_38_18 (
    .O(x38_y18),
    .I0(x36_y14),
    .I1(x35_y15),
    .I2(x35_y21),
    .I3(x35_y15)
);

(* keep, dont_touch *)
(* LOC = "X39/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000010110101)
) lut_39_18 (
    .O(x39_y18),
    .I0(1'b0),
    .I1(x37_y14),
    .I2(1'b0),
    .I3(x37_y21)
);

(* keep, dont_touch *)
(* LOC = "X40/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100101110111)
) lut_40_18 (
    .O(x40_y18),
    .I0(1'b0),
    .I1(x38_y15),
    .I2(1'b0),
    .I3(x38_y23)
);

(* keep, dont_touch *)
(* LOC = "X41/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111001010110)
) lut_41_18 (
    .O(x41_y18),
    .I0(x39_y15),
    .I1(1'b0),
    .I2(x39_y18),
    .I3(x39_y18)
);

(* keep, dont_touch *)
(* LOC = "X42/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010110101001)
) lut_42_18 (
    .O(x42_y18),
    .I0(x40_y13),
    .I1(x40_y17),
    .I2(1'b0),
    .I3(x39_y19)
);

(* keep, dont_touch *)
(* LOC = "X43/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110011001101)
) lut_43_18 (
    .O(x43_y18),
    .I0(x41_y19),
    .I1(x40_y21),
    .I2(x40_y22),
    .I3(x40_y17)
);

(* keep, dont_touch *)
(* LOC = "X44/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000111001001)
) lut_44_18 (
    .O(x44_y18),
    .I0(1'b0),
    .I1(x42_y23),
    .I2(1'b0),
    .I3(x42_y16)
);

(* keep, dont_touch *)
(* LOC = "X45/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100100100010)
) lut_45_18 (
    .O(x45_y18),
    .I0(x42_y16),
    .I1(x43_y13),
    .I2(x43_y22),
    .I3(x43_y21)
);

(* keep, dont_touch *)
(* LOC = "X46/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010010110111)
) lut_46_18 (
    .O(x46_y18),
    .I0(x44_y23),
    .I1(x43_y19),
    .I2(x43_y18),
    .I3(x43_y21)
);

(* keep, dont_touch *)
(* LOC = "X47/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011001111100)
) lut_47_18 (
    .O(x47_y18),
    .I0(x44_y17),
    .I1(1'b0),
    .I2(x44_y16),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X48/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011100110001)
) lut_48_18 (
    .O(x48_y18),
    .I0(1'b0),
    .I1(x45_y14),
    .I2(x46_y19),
    .I3(x46_y21)
);

(* keep, dont_touch *)
(* LOC = "X49/Y18" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111100100010)
) lut_49_18 (
    .O(x49_y18),
    .I0(x47_y17),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x47_y21)
);

(* keep, dont_touch *)
(* LOC = "X0/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101101111101)
) lut_0_19 (
    .O(x0_y19),
    .I0(in8),
    .I1(in4),
    .I2(in5),
    .I3(in3)
);

(* keep, dont_touch *)
(* LOC = "X1/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100001000100)
) lut_1_19 (
    .O(x1_y19),
    .I0(in0),
    .I1(in2),
    .I2(in9),
    .I3(in8)
);

(* keep, dont_touch *)
(* LOC = "X2/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101100000100)
) lut_2_19 (
    .O(x2_y19),
    .I0(in1),
    .I1(in7),
    .I2(1'b0),
    .I3(in6)
);

(* keep, dont_touch *)
(* LOC = "X3/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110100011101)
) lut_3_19 (
    .O(x3_y19),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x1_y20),
    .I3(x1_y21)
);

(* keep, dont_touch *)
(* LOC = "X4/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001111100001)
) lut_4_19 (
    .O(x4_y19),
    .I0(x2_y20),
    .I1(x1_y24),
    .I2(1'b0),
    .I3(x2_y24)
);

(* keep, dont_touch *)
(* LOC = "X5/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111000111011)
) lut_5_19 (
    .O(x5_y19),
    .I0(1'b0),
    .I1(x3_y19),
    .I2(x2_y17),
    .I3(x3_y23)
);

(* keep, dont_touch *)
(* LOC = "X6/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101111100111)
) lut_6_19 (
    .O(x6_y19),
    .I0(x4_y21),
    .I1(1'b0),
    .I2(x4_y23),
    .I3(x4_y20)
);

(* keep, dont_touch *)
(* LOC = "X7/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011010010011)
) lut_7_19 (
    .O(x7_y19),
    .I0(x5_y15),
    .I1(x5_y17),
    .I2(x5_y21),
    .I3(x5_y21)
);

(* keep, dont_touch *)
(* LOC = "X8/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001001101110)
) lut_8_19 (
    .O(x8_y19),
    .I0(x6_y24),
    .I1(x6_y17),
    .I2(1'b0),
    .I3(x6_y21)
);

(* keep, dont_touch *)
(* LOC = "X9/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000110011101)
) lut_9_19 (
    .O(x9_y19),
    .I0(x6_y20),
    .I1(x7_y22),
    .I2(1'b0),
    .I3(x6_y21)
);

(* keep, dont_touch *)
(* LOC = "X10/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010000000100)
) lut_10_19 (
    .O(x10_y19),
    .I0(1'b0),
    .I1(x8_y24),
    .I2(x7_y21),
    .I3(x8_y24)
);

(* keep, dont_touch *)
(* LOC = "X11/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110011001111)
) lut_11_19 (
    .O(x11_y19),
    .I0(x8_y20),
    .I1(x9_y19),
    .I2(x9_y16),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X12/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000011110110)
) lut_12_19 (
    .O(x12_y19),
    .I0(x10_y14),
    .I1(1'b0),
    .I2(x9_y23),
    .I3(x10_y17)
);

(* keep, dont_touch *)
(* LOC = "X13/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111001000111)
) lut_13_19 (
    .O(x13_y19),
    .I0(x10_y15),
    .I1(x11_y20),
    .I2(1'b0),
    .I3(x11_y18)
);

(* keep, dont_touch *)
(* LOC = "X14/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100111111001)
) lut_14_19 (
    .O(x14_y19),
    .I0(x11_y23),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x11_y22)
);

(* keep, dont_touch *)
(* LOC = "X15/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100011111000)
) lut_15_19 (
    .O(x15_y19),
    .I0(x13_y23),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x13_y24)
);

(* keep, dont_touch *)
(* LOC = "X16/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000011000100)
) lut_16_19 (
    .O(x16_y19),
    .I0(x14_y20),
    .I1(x13_y15),
    .I2(x13_y18),
    .I3(x13_y17)
);

(* keep, dont_touch *)
(* LOC = "X17/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111100010001)
) lut_17_19 (
    .O(x17_y19),
    .I0(x14_y18),
    .I1(x15_y21),
    .I2(1'b0),
    .I3(x15_y15)
);

(* keep, dont_touch *)
(* LOC = "X18/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111011100010)
) lut_18_19 (
    .O(x18_y19),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x16_y24),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X19/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010001000101)
) lut_19_19 (
    .O(x19_y19),
    .I0(x16_y18),
    .I1(x17_y20),
    .I2(x17_y17),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X20/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110111011001)
) lut_20_19 (
    .O(x20_y19),
    .I0(x17_y24),
    .I1(1'b0),
    .I2(x17_y21),
    .I3(x18_y18)
);

(* keep, dont_touch *)
(* LOC = "X21/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001010100001)
) lut_21_19 (
    .O(x21_y19),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x19_y21),
    .I3(x19_y21)
);

(* keep, dont_touch *)
(* LOC = "X22/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001011100000)
) lut_22_19 (
    .O(x22_y19),
    .I0(x20_y15),
    .I1(x19_y17),
    .I2(1'b0),
    .I3(x20_y16)
);

(* keep, dont_touch *)
(* LOC = "X23/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100010000110)
) lut_23_19 (
    .O(x23_y19),
    .I0(x21_y18),
    .I1(x20_y23),
    .I2(x20_y23),
    .I3(x20_y15)
);

(* keep, dont_touch *)
(* LOC = "X24/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100001100101)
) lut_24_19 (
    .O(x24_y19),
    .I0(1'b0),
    .I1(x22_y16),
    .I2(x22_y24),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X25/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110001010001)
) lut_25_19 (
    .O(x25_y19),
    .I0(x23_y22),
    .I1(x22_y14),
    .I2(1'b0),
    .I3(x23_y20)
);

(* keep, dont_touch *)
(* LOC = "X26/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100100000100)
) lut_26_19 (
    .O(x26_y19),
    .I0(x23_y24),
    .I1(1'b0),
    .I2(x23_y15),
    .I3(x23_y21)
);

(* keep, dont_touch *)
(* LOC = "X27/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110000011010)
) lut_27_19 (
    .O(x27_y19),
    .I0(x25_y23),
    .I1(x24_y22),
    .I2(x24_y18),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X28/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101110100110)
) lut_28_19 (
    .O(x28_y19),
    .I0(x25_y19),
    .I1(1'b0),
    .I2(x26_y24),
    .I3(x25_y21)
);

(* keep, dont_touch *)
(* LOC = "X29/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110010111110)
) lut_29_19 (
    .O(x29_y19),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x26_y16),
    .I3(x27_y23)
);

(* keep, dont_touch *)
(* LOC = "X30/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000000110101)
) lut_30_19 (
    .O(x30_y19),
    .I0(x27_y23),
    .I1(x28_y17),
    .I2(x28_y19),
    .I3(x27_y20)
);

(* keep, dont_touch *)
(* LOC = "X31/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101001000111)
) lut_31_19 (
    .O(x31_y19),
    .I0(x29_y20),
    .I1(x29_y18),
    .I2(x29_y15),
    .I3(x29_y15)
);

(* keep, dont_touch *)
(* LOC = "X32/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011100011100)
) lut_32_19 (
    .O(x32_y19),
    .I0(x29_y20),
    .I1(x29_y14),
    .I2(x30_y19),
    .I3(x30_y21)
);

(* keep, dont_touch *)
(* LOC = "X33/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011101101100)
) lut_33_19 (
    .O(x33_y19),
    .I0(x31_y18),
    .I1(1'b0),
    .I2(x31_y15),
    .I3(x31_y16)
);

(* keep, dont_touch *)
(* LOC = "X34/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111000001011)
) lut_34_19 (
    .O(x34_y19),
    .I0(x31_y14),
    .I1(1'b0),
    .I2(x31_y21),
    .I3(x32_y15)
);

(* keep, dont_touch *)
(* LOC = "X35/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110100110101)
) lut_35_19 (
    .O(x35_y19),
    .I0(x32_y24),
    .I1(1'b0),
    .I2(x32_y16),
    .I3(x33_y18)
);

(* keep, dont_touch *)
(* LOC = "X36/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000100100010)
) lut_36_19 (
    .O(x36_y19),
    .I0(x33_y15),
    .I1(x33_y21),
    .I2(x34_y22),
    .I3(x34_y21)
);

(* keep, dont_touch *)
(* LOC = "X37/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111110011011)
) lut_37_19 (
    .O(x37_y19),
    .I0(x35_y16),
    .I1(x35_y21),
    .I2(x35_y18),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X38/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110010010101)
) lut_38_19 (
    .O(x38_y19),
    .I0(x35_y16),
    .I1(1'b0),
    .I2(x36_y20),
    .I3(x35_y21)
);

(* keep, dont_touch *)
(* LOC = "X39/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100101110100)
) lut_39_19 (
    .O(x39_y19),
    .I0(x37_y16),
    .I1(x37_y14),
    .I2(1'b0),
    .I3(x36_y20)
);

(* keep, dont_touch *)
(* LOC = "X40/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011100111011)
) lut_40_19 (
    .O(x40_y19),
    .I0(1'b0),
    .I1(x38_y18),
    .I2(x38_y17),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X41/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000000111011)
) lut_41_19 (
    .O(x41_y19),
    .I0(1'b0),
    .I1(x38_y21),
    .I2(1'b0),
    .I3(x38_y22)
);

(* keep, dont_touch *)
(* LOC = "X42/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110111001100)
) lut_42_19 (
    .O(x42_y19),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x40_y21)
);

(* keep, dont_touch *)
(* LOC = "X43/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011111110010)
) lut_43_19 (
    .O(x43_y19),
    .I0(1'b0),
    .I1(x41_y16),
    .I2(x40_y24),
    .I3(x40_y23)
);

(* keep, dont_touch *)
(* LOC = "X44/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011111010000)
) lut_44_19 (
    .O(x44_y19),
    .I0(x41_y19),
    .I1(x41_y21),
    .I2(x42_y16),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X45/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110010001010)
) lut_45_19 (
    .O(x45_y19),
    .I0(x43_y24),
    .I1(x42_y21),
    .I2(x42_y16),
    .I3(x42_y23)
);

(* keep, dont_touch *)
(* LOC = "X46/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010111010011)
) lut_46_19 (
    .O(x46_y19),
    .I0(x44_y19),
    .I1(x44_y22),
    .I2(x44_y22),
    .I3(x44_y23)
);

(* keep, dont_touch *)
(* LOC = "X47/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001110100001)
) lut_47_19 (
    .O(x47_y19),
    .I0(x44_y19),
    .I1(x44_y22),
    .I2(x45_y16),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X48/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101111001001)
) lut_48_19 (
    .O(x48_y19),
    .I0(x46_y21),
    .I1(1'b0),
    .I2(x45_y24),
    .I3(x45_y16)
);

(* keep, dont_touch *)
(* LOC = "X49/Y19" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110010011000)
) lut_49_19 (
    .O(x49_y19),
    .I0(x46_y22),
    .I1(x46_y16),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X0/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000010000001)
) lut_0_20 (
    .O(x0_y20),
    .I0(in5),
    .I1(in5),
    .I2(in0),
    .I3(in4)
);

(* keep, dont_touch *)
(* LOC = "X1/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110101111011)
) lut_1_20 (
    .O(x1_y20),
    .I0(in0),
    .I1(in5),
    .I2(in6),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X2/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111111011101)
) lut_2_20 (
    .O(x2_y20),
    .I0(in2),
    .I1(in0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X3/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011001110111)
) lut_3_20 (
    .O(x3_y20),
    .I0(x1_y24),
    .I1(1'b0),
    .I2(in5),
    .I3(in6)
);

(* keep, dont_touch *)
(* LOC = "X4/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100011110001)
) lut_4_20 (
    .O(x4_y20),
    .I0(1'b0),
    .I1(x1_y15),
    .I2(1'b0),
    .I3(x1_y19)
);

(* keep, dont_touch *)
(* LOC = "X5/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001110010111)
) lut_5_20 (
    .O(x5_y20),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x3_y15),
    .I3(x3_y23)
);

(* keep, dont_touch *)
(* LOC = "X6/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110000101111)
) lut_6_20 (
    .O(x6_y20),
    .I0(x4_y23),
    .I1(x3_y25),
    .I2(x3_y16),
    .I3(x4_y15)
);

(* keep, dont_touch *)
(* LOC = "X7/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011101101010)
) lut_7_20 (
    .O(x7_y20),
    .I0(x4_y16),
    .I1(x5_y20),
    .I2(x5_y22),
    .I3(x5_y20)
);

(* keep, dont_touch *)
(* LOC = "X8/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010001011001)
) lut_8_20 (
    .O(x8_y20),
    .I0(x5_y19),
    .I1(x6_y17),
    .I2(x6_y24),
    .I3(x6_y21)
);

(* keep, dont_touch *)
(* LOC = "X9/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111001101101)
) lut_9_20 (
    .O(x9_y20),
    .I0(x7_y15),
    .I1(x7_y19),
    .I2(x6_y24),
    .I3(x6_y21)
);

(* keep, dont_touch *)
(* LOC = "X10/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101010001001)
) lut_10_20 (
    .O(x10_y20),
    .I0(x8_y17),
    .I1(x8_y22),
    .I2(x8_y24),
    .I3(x7_y15)
);

(* keep, dont_touch *)
(* LOC = "X11/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111100101001)
) lut_11_20 (
    .O(x11_y20),
    .I0(x8_y23),
    .I1(x8_y19),
    .I2(x8_y17),
    .I3(x9_y17)
);

(* keep, dont_touch *)
(* LOC = "X12/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101001101011)
) lut_12_20 (
    .O(x12_y20),
    .I0(1'b0),
    .I1(x10_y22),
    .I2(1'b0),
    .I3(x9_y16)
);

(* keep, dont_touch *)
(* LOC = "X13/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010011101010)
) lut_13_20 (
    .O(x13_y20),
    .I0(x10_y22),
    .I1(x10_y20),
    .I2(1'b0),
    .I3(x10_y22)
);

(* keep, dont_touch *)
(* LOC = "X14/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011111110101)
) lut_14_20 (
    .O(x14_y20),
    .I0(x11_y15),
    .I1(x12_y19),
    .I2(1'b0),
    .I3(x12_y21)
);

(* keep, dont_touch *)
(* LOC = "X15/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101101011010)
) lut_15_20 (
    .O(x15_y20),
    .I0(1'b0),
    .I1(x13_y15),
    .I2(x13_y25),
    .I3(x13_y16)
);

(* keep, dont_touch *)
(* LOC = "X16/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100000101101)
) lut_16_20 (
    .O(x16_y20),
    .I0(1'b0),
    .I1(x14_y15),
    .I2(x13_y16),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X17/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010010000010)
) lut_17_20 (
    .O(x17_y20),
    .I0(x14_y17),
    .I1(x14_y24),
    .I2(x14_y20),
    .I3(x14_y16)
);

(* keep, dont_touch *)
(* LOC = "X18/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011010000011)
) lut_18_20 (
    .O(x18_y20),
    .I0(1'b0),
    .I1(x16_y21),
    .I2(x15_y16),
    .I3(x16_y17)
);

(* keep, dont_touch *)
(* LOC = "X19/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100000001000)
) lut_19_20 (
    .O(x19_y20),
    .I0(x16_y21),
    .I1(x16_y25),
    .I2(x17_y19),
    .I3(x17_y24)
);

(* keep, dont_touch *)
(* LOC = "X20/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110110010100)
) lut_20_20 (
    .O(x20_y20),
    .I0(x17_y24),
    .I1(1'b0),
    .I2(x17_y21),
    .I3(x18_y19)
);

(* keep, dont_touch *)
(* LOC = "X21/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010000000101)
) lut_21_20 (
    .O(x21_y20),
    .I0(x19_y19),
    .I1(x19_y25),
    .I2(x18_y21),
    .I3(x19_y20)
);

(* keep, dont_touch *)
(* LOC = "X22/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101001100001)
) lut_22_20 (
    .O(x22_y20),
    .I0(x20_y15),
    .I1(x20_y24),
    .I2(x20_y23),
    .I3(x20_y22)
);

(* keep, dont_touch *)
(* LOC = "X23/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010110110010)
) lut_23_20 (
    .O(x23_y20),
    .I0(x20_y24),
    .I1(x21_y23),
    .I2(x20_y18),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X24/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100001011001)
) lut_24_20 (
    .O(x24_y20),
    .I0(x21_y15),
    .I1(x22_y16),
    .I2(x22_y15),
    .I3(x21_y19)
);

(* keep, dont_touch *)
(* LOC = "X25/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001111100000)
) lut_25_20 (
    .O(x25_y20),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x22_y15),
    .I3(x23_y24)
);

(* keep, dont_touch *)
(* LOC = "X26/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010010101101)
) lut_26_20 (
    .O(x26_y20),
    .I0(x23_y18),
    .I1(x24_y18),
    .I2(x24_y20),
    .I3(x23_y23)
);

(* keep, dont_touch *)
(* LOC = "X27/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011111100000)
) lut_27_20 (
    .O(x27_y20),
    .I0(x24_y21),
    .I1(x25_y21),
    .I2(x25_y22),
    .I3(x25_y21)
);

(* keep, dont_touch *)
(* LOC = "X28/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011100100101)
) lut_28_20 (
    .O(x28_y20),
    .I0(1'b0),
    .I1(x26_y19),
    .I2(x26_y15),
    .I3(x25_y18)
);

(* keep, dont_touch *)
(* LOC = "X29/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101101010010)
) lut_29_20 (
    .O(x29_y20),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x26_y23),
    .I3(x26_y15)
);

(* keep, dont_touch *)
(* LOC = "X30/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110011111110)
) lut_30_20 (
    .O(x30_y20),
    .I0(1'b0),
    .I1(x27_y17),
    .I2(x27_y23),
    .I3(x27_y23)
);

(* keep, dont_touch *)
(* LOC = "X31/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001010001110)
) lut_31_20 (
    .O(x31_y20),
    .I0(x29_y22),
    .I1(x28_y24),
    .I2(x28_y20),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X32/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100110111100)
) lut_32_20 (
    .O(x32_y20),
    .I0(x29_y17),
    .I1(1'b0),
    .I2(x29_y19),
    .I3(x30_y20)
);

(* keep, dont_touch *)
(* LOC = "X33/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010111101100)
) lut_33_20 (
    .O(x33_y20),
    .I0(1'b0),
    .I1(x31_y16),
    .I2(x30_y17),
    .I3(x30_y20)
);

(* keep, dont_touch *)
(* LOC = "X34/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101001110111)
) lut_34_20 (
    .O(x34_y20),
    .I0(x31_y24),
    .I1(x32_y21),
    .I2(1'b0),
    .I3(x32_y16)
);

(* keep, dont_touch *)
(* LOC = "X35/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111001001000)
) lut_35_20 (
    .O(x35_y20),
    .I0(x33_y16),
    .I1(x33_y19),
    .I2(1'b0),
    .I3(x32_y23)
);

(* keep, dont_touch *)
(* LOC = "X36/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101000100000)
) lut_36_20 (
    .O(x36_y20),
    .I0(x34_y15),
    .I1(x33_y15),
    .I2(1'b0),
    .I3(x33_y24)
);

(* keep, dont_touch *)
(* LOC = "X37/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110111100111)
) lut_37_20 (
    .O(x37_y20),
    .I0(x35_y23),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x35_y21)
);

(* keep, dont_touch *)
(* LOC = "X38/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011100110110)
) lut_38_20 (
    .O(x38_y20),
    .I0(1'b0),
    .I1(x35_y21),
    .I2(x35_y24),
    .I3(x36_y20)
);

(* keep, dont_touch *)
(* LOC = "X39/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011001011110)
) lut_39_20 (
    .O(x39_y20),
    .I0(x36_y25),
    .I1(1'b0),
    .I2(x37_y24),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X40/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011110111101)
) lut_40_20 (
    .O(x40_y20),
    .I0(x37_y20),
    .I1(x38_y25),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X41/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010000001011)
) lut_41_20 (
    .O(x41_y20),
    .I0(x38_y23),
    .I1(1'b0),
    .I2(x38_y19),
    .I3(x39_y24)
);

(* keep, dont_touch *)
(* LOC = "X42/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010110001110)
) lut_42_20 (
    .O(x42_y20),
    .I0(x40_y19),
    .I1(1'b0),
    .I2(x40_y24),
    .I3(x40_y18)
);

(* keep, dont_touch *)
(* LOC = "X43/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001000000010)
) lut_43_20 (
    .O(x43_y20),
    .I0(1'b0),
    .I1(x41_y15),
    .I2(1'b0),
    .I3(x40_y21)
);

(* keep, dont_touch *)
(* LOC = "X44/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101011011011)
) lut_44_20 (
    .O(x44_y20),
    .I0(x41_y18),
    .I1(x42_y21),
    .I2(x42_y15),
    .I3(x41_y22)
);

(* keep, dont_touch *)
(* LOC = "X45/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011011010110)
) lut_45_20 (
    .O(x45_y20),
    .I0(x43_y19),
    .I1(1'b0),
    .I2(x43_y24),
    .I3(x42_y25)
);

(* keep, dont_touch *)
(* LOC = "X46/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111001101101)
) lut_46_20 (
    .O(x46_y20),
    .I0(x43_y22),
    .I1(1'b0),
    .I2(x44_y22),
    .I3(x44_y21)
);

(* keep, dont_touch *)
(* LOC = "X47/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111101001000)
) lut_47_20 (
    .O(x47_y20),
    .I0(1'b0),
    .I1(x44_y19),
    .I2(x44_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X48/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001101010111)
) lut_48_20 (
    .O(x48_y20),
    .I0(x46_y21),
    .I1(x46_y24),
    .I2(x46_y15),
    .I3(x45_y23)
);

(* keep, dont_touch *)
(* LOC = "X49/Y20" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111011110101)
) lut_49_20 (
    .O(x49_y20),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x47_y17),
    .I3(x46_y17)
);

(* keep, dont_touch *)
(* LOC = "X0/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010010001101)
) lut_0_21 (
    .O(x0_y21),
    .I0(in2),
    .I1(in6),
    .I2(1'b0),
    .I3(in8)
);

(* keep, dont_touch *)
(* LOC = "X1/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001011001100)
) lut_1_21 (
    .O(x1_y21),
    .I0(in2),
    .I1(1'b0),
    .I2(in3),
    .I3(in5)
);

(* keep, dont_touch *)
(* LOC = "X2/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100111000100)
) lut_2_21 (
    .O(x2_y21),
    .I0(in4),
    .I1(in3),
    .I2(in5),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X3/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010101110101)
) lut_3_21 (
    .O(x3_y21),
    .I0(1'b0),
    .I1(x1_y26),
    .I2(x1_y18),
    .I3(x1_y26)
);

(* keep, dont_touch *)
(* LOC = "X4/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110100100100)
) lut_4_21 (
    .O(x4_y21),
    .I0(1'b0),
    .I1(x1_y26),
    .I2(x2_y17),
    .I3(x2_y26)
);

(* keep, dont_touch *)
(* LOC = "X5/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011011100001)
) lut_5_21 (
    .O(x5_y21),
    .I0(x3_y25),
    .I1(x3_y20),
    .I2(x2_y19),
    .I3(x2_y17)
);

(* keep, dont_touch *)
(* LOC = "X6/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100101101010)
) lut_6_21 (
    .O(x6_y21),
    .I0(1'b0),
    .I1(x3_y26),
    .I2(x4_y20),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X7/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011100101000)
) lut_7_21 (
    .O(x7_y21),
    .I0(x5_y19),
    .I1(x5_y19),
    .I2(x5_y23),
    .I3(x5_y26)
);

(* keep, dont_touch *)
(* LOC = "X8/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110111110111)
) lut_8_21 (
    .O(x8_y21),
    .I0(x5_y18),
    .I1(x6_y25),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X9/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110000111000)
) lut_9_21 (
    .O(x9_y21),
    .I0(x6_y23),
    .I1(x7_y20),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X10/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110111110000)
) lut_10_21 (
    .O(x10_y21),
    .I0(x7_y19),
    .I1(x8_y24),
    .I2(x8_y22),
    .I3(x7_y16)
);

(* keep, dont_touch *)
(* LOC = "X11/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101001000111)
) lut_11_21 (
    .O(x11_y21),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x9_y23),
    .I3(x9_y20)
);

(* keep, dont_touch *)
(* LOC = "X12/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100110110001)
) lut_12_21 (
    .O(x12_y21),
    .I0(x10_y18),
    .I1(x10_y19),
    .I2(x10_y22),
    .I3(x10_y22)
);

(* keep, dont_touch *)
(* LOC = "X13/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110111000010)
) lut_13_21 (
    .O(x13_y21),
    .I0(x10_y17),
    .I1(x11_y19),
    .I2(x10_y16),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X14/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111111000001)
) lut_14_21 (
    .O(x14_y21),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x12_y26),
    .I3(x12_y19)
);

(* keep, dont_touch *)
(* LOC = "X15/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000010001110)
) lut_15_21 (
    .O(x15_y21),
    .I0(1'b0),
    .I1(x12_y17),
    .I2(x13_y17),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X16/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010010101101)
) lut_16_21 (
    .O(x16_y21),
    .I0(x14_y16),
    .I1(x13_y25),
    .I2(1'b0),
    .I3(x13_y24)
);

(* keep, dont_touch *)
(* LOC = "X17/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110110000100)
) lut_17_21 (
    .O(x17_y21),
    .I0(x14_y21),
    .I1(x15_y20),
    .I2(x15_y16),
    .I3(x15_y17)
);

(* keep, dont_touch *)
(* LOC = "X18/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010101100111)
) lut_18_21 (
    .O(x18_y21),
    .I0(x15_y24),
    .I1(x15_y24),
    .I2(x15_y21),
    .I3(x15_y19)
);

(* keep, dont_touch *)
(* LOC = "X19/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111010001010)
) lut_19_21 (
    .O(x19_y21),
    .I0(1'b0),
    .I1(x17_y17),
    .I2(1'b0),
    .I3(x16_y26)
);

(* keep, dont_touch *)
(* LOC = "X20/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001111010000)
) lut_20_21 (
    .O(x20_y21),
    .I0(x18_y25),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x18_y22)
);

(* keep, dont_touch *)
(* LOC = "X21/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011101100000)
) lut_21_21 (
    .O(x21_y21),
    .I0(x18_y23),
    .I1(1'b0),
    .I2(x18_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X22/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100100000000)
) lut_22_21 (
    .O(x22_y21),
    .I0(x19_y21),
    .I1(x20_y18),
    .I2(x20_y23),
    .I3(x19_y23)
);

(* keep, dont_touch *)
(* LOC = "X23/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001101011001)
) lut_23_21 (
    .O(x23_y21),
    .I0(x20_y17),
    .I1(x21_y17),
    .I2(x21_y23),
    .I3(x20_y24)
);

(* keep, dont_touch *)
(* LOC = "X24/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011111010010)
) lut_24_21 (
    .O(x24_y21),
    .I0(1'b0),
    .I1(x22_y21),
    .I2(x22_y17),
    .I3(x22_y24)
);

(* keep, dont_touch *)
(* LOC = "X25/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111110110110)
) lut_25_21 (
    .O(x25_y21),
    .I0(x22_y24),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x22_y26)
);

(* keep, dont_touch *)
(* LOC = "X26/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101101011100)
) lut_26_21 (
    .O(x26_y21),
    .I0(x24_y24),
    .I1(x23_y24),
    .I2(x23_y24),
    .I3(x23_y25)
);

(* keep, dont_touch *)
(* LOC = "X27/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000000011000)
) lut_27_21 (
    .O(x27_y21),
    .I0(x25_y17),
    .I1(x24_y16),
    .I2(x25_y19),
    .I3(x25_y18)
);

(* keep, dont_touch *)
(* LOC = "X28/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001010100110)
) lut_28_21 (
    .O(x28_y21),
    .I0(x26_y21),
    .I1(1'b0),
    .I2(x25_y17),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X29/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000101101110)
) lut_29_21 (
    .O(x29_y21),
    .I0(x27_y24),
    .I1(x26_y24),
    .I2(1'b0),
    .I3(x27_y20)
);

(* keep, dont_touch *)
(* LOC = "X30/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101111000100)
) lut_30_21 (
    .O(x30_y21),
    .I0(x28_y16),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x28_y17)
);

(* keep, dont_touch *)
(* LOC = "X31/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010010001010)
) lut_31_21 (
    .O(x31_y21),
    .I0(x28_y22),
    .I1(1'b0),
    .I2(x29_y16),
    .I3(x28_y23)
);

(* keep, dont_touch *)
(* LOC = "X32/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100100110000)
) lut_32_21 (
    .O(x32_y21),
    .I0(x30_y19),
    .I1(1'b0),
    .I2(x29_y19),
    .I3(x29_y21)
);

(* keep, dont_touch *)
(* LOC = "X33/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100101010111)
) lut_33_21 (
    .O(x33_y21),
    .I0(x30_y22),
    .I1(1'b0),
    .I2(x30_y20),
    .I3(x31_y26)
);

(* keep, dont_touch *)
(* LOC = "X34/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101010110101)
) lut_34_21 (
    .O(x34_y21),
    .I0(x32_y26),
    .I1(x32_y22),
    .I2(x32_y25),
    .I3(x31_y25)
);

(* keep, dont_touch *)
(* LOC = "X35/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011101001001)
) lut_35_21 (
    .O(x35_y21),
    .I0(x32_y22),
    .I1(x32_y16),
    .I2(x32_y17),
    .I3(x32_y23)
);

(* keep, dont_touch *)
(* LOC = "X36/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001010000101)
) lut_36_21 (
    .O(x36_y21),
    .I0(x33_y25),
    .I1(x34_y21),
    .I2(1'b0),
    .I3(x33_y21)
);

(* keep, dont_touch *)
(* LOC = "X37/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111001110101)
) lut_37_21 (
    .O(x37_y21),
    .I0(x34_y24),
    .I1(x34_y17),
    .I2(x35_y18),
    .I3(x34_y25)
);

(* keep, dont_touch *)
(* LOC = "X38/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100001000101)
) lut_38_21 (
    .O(x38_y21),
    .I0(x36_y16),
    .I1(1'b0),
    .I2(x35_y23),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X39/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101100010110)
) lut_39_21 (
    .O(x39_y21),
    .I0(x36_y21),
    .I1(x36_y23),
    .I2(x37_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X40/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010110110101)
) lut_40_21 (
    .O(x40_y21),
    .I0(x37_y26),
    .I1(x38_y26),
    .I2(x38_y18),
    .I3(x37_y20)
);

(* keep, dont_touch *)
(* LOC = "X41/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001101101001)
) lut_41_21 (
    .O(x41_y21),
    .I0(x38_y22),
    .I1(x39_y19),
    .I2(x39_y18),
    .I3(x39_y16)
);

(* keep, dont_touch *)
(* LOC = "X42/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101100000111)
) lut_42_21 (
    .O(x42_y21),
    .I0(1'b0),
    .I1(x40_y25),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X43/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011011001111)
) lut_43_21 (
    .O(x43_y21),
    .I0(x40_y17),
    .I1(x40_y18),
    .I2(x40_y20),
    .I3(x40_y24)
);

(* keep, dont_touch *)
(* LOC = "X44/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000101110101)
) lut_44_21 (
    .O(x44_y21),
    .I0(x42_y17),
    .I1(x41_y26),
    .I2(x41_y24),
    .I3(x41_y25)
);

(* keep, dont_touch *)
(* LOC = "X45/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111000001010)
) lut_45_21 (
    .O(x45_y21),
    .I0(x43_y26),
    .I1(x42_y23),
    .I2(x42_y18),
    .I3(x43_y25)
);

(* keep, dont_touch *)
(* LOC = "X46/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010011000011)
) lut_46_21 (
    .O(x46_y21),
    .I0(x44_y24),
    .I1(1'b0),
    .I2(x43_y17),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X47/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101001110001)
) lut_47_21 (
    .O(x47_y21),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x45_y17),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X48/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001011010110)
) lut_48_21 (
    .O(x48_y21),
    .I0(x46_y20),
    .I1(1'b0),
    .I2(x45_y23),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X49/Y21" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001110100000)
) lut_49_21 (
    .O(x49_y21),
    .I0(x46_y23),
    .I1(x47_y26),
    .I2(x46_y21),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X0/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000111110110)
) lut_0_22 (
    .O(x0_y22),
    .I0(1'b0),
    .I1(in8),
    .I2(in2),
    .I3(in4)
);

(* keep, dont_touch *)
(* LOC = "X1/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101000100100)
) lut_1_22 (
    .O(x1_y22),
    .I0(in9),
    .I1(1'b0),
    .I2(in7),
    .I3(in1)
);

(* keep, dont_touch *)
(* LOC = "X2/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110101000100)
) lut_2_22 (
    .O(x2_y22),
    .I0(in7),
    .I1(in5),
    .I2(in0),
    .I3(in6)
);

(* keep, dont_touch *)
(* LOC = "X3/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010101100000)
) lut_3_22 (
    .O(x3_y22),
    .I0(x1_y24),
    .I1(1'b0),
    .I2(in0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X4/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110101011010)
) lut_4_22 (
    .O(x4_y22),
    .I0(x1_y17),
    .I1(x1_y21),
    .I2(x2_y23),
    .I3(x2_y18)
);

(* keep, dont_touch *)
(* LOC = "X5/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111100100110)
) lut_5_22 (
    .O(x5_y22),
    .I0(1'b0),
    .I1(x3_y23),
    .I2(x3_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X6/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101100011101)
) lut_6_22 (
    .O(x6_y22),
    .I0(x3_y20),
    .I1(x3_y23),
    .I2(x3_y17),
    .I3(x3_y26)
);

(* keep, dont_touch *)
(* LOC = "X7/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100111001111)
) lut_7_22 (
    .O(x7_y22),
    .I0(1'b0),
    .I1(x5_y27),
    .I2(x5_y22),
    .I3(x4_y19)
);

(* keep, dont_touch *)
(* LOC = "X8/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100101001111)
) lut_8_22 (
    .O(x8_y22),
    .I0(x6_y20),
    .I1(x6_y22),
    .I2(x5_y27),
    .I3(x5_y21)
);

(* keep, dont_touch *)
(* LOC = "X9/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000001011000)
) lut_9_22 (
    .O(x9_y22),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x5_y27),
    .I3(x5_y21)
);

(* keep, dont_touch *)
(* LOC = "X10/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111111111111)
) lut_10_22 (
    .O(x10_y22),
    .I0(1'b0),
    .I1(x8_y22),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X11/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010010010001)
) lut_11_22 (
    .O(x11_y22),
    .I0(x9_y23),
    .I1(1'b0),
    .I2(x9_y21),
    .I3(x8_y18)
);

(* keep, dont_touch *)
(* LOC = "X12/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011100011100)
) lut_12_22 (
    .O(x12_y22),
    .I0(x9_y27),
    .I1(x9_y25),
    .I2(1'b0),
    .I3(x10_y27)
);

(* keep, dont_touch *)
(* LOC = "X13/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100100100101)
) lut_13_22 (
    .O(x13_y22),
    .I0(x10_y23),
    .I1(1'b0),
    .I2(x11_y23),
    .I3(x11_y26)
);

(* keep, dont_touch *)
(* LOC = "X14/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010101100011)
) lut_14_22 (
    .O(x14_y22),
    .I0(x12_y24),
    .I1(x11_y22),
    .I2(x11_y23),
    .I3(x11_y17)
);

(* keep, dont_touch *)
(* LOC = "X15/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010001110100)
) lut_15_22 (
    .O(x15_y22),
    .I0(x13_y24),
    .I1(x12_y21),
    .I2(1'b0),
    .I3(x13_y18)
);

(* keep, dont_touch *)
(* LOC = "X16/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101110100001)
) lut_16_22 (
    .O(x16_y22),
    .I0(x14_y21),
    .I1(x13_y19),
    .I2(x14_y24),
    .I3(x13_y22)
);

(* keep, dont_touch *)
(* LOC = "X17/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111100100011)
) lut_17_22 (
    .O(x17_y22),
    .I0(x15_y25),
    .I1(x15_y27),
    .I2(x15_y25),
    .I3(x14_y27)
);

(* keep, dont_touch *)
(* LOC = "X18/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100010011111)
) lut_18_22 (
    .O(x18_y22),
    .I0(x16_y19),
    .I1(x16_y19),
    .I2(x16_y25),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X19/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100000111111)
) lut_19_22 (
    .O(x19_y22),
    .I0(1'b0),
    .I1(x17_y27),
    .I2(x17_y27),
    .I3(x16_y23)
);

(* keep, dont_touch *)
(* LOC = "X20/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001000000011)
) lut_20_22 (
    .O(x20_y22),
    .I0(x17_y22),
    .I1(x17_y18),
    .I2(x17_y26),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X21/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101010100010)
) lut_21_22 (
    .O(x21_y22),
    .I0(x18_y17),
    .I1(x19_y18),
    .I2(x18_y20),
    .I3(x19_y21)
);

(* keep, dont_touch *)
(* LOC = "X22/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101000101000)
) lut_22_22 (
    .O(x22_y22),
    .I0(x19_y21),
    .I1(x19_y25),
    .I2(x20_y21),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X23/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000101110101)
) lut_23_22 (
    .O(x23_y22),
    .I0(x20_y27),
    .I1(x20_y27),
    .I2(x20_y19),
    .I3(x21_y27)
);

(* keep, dont_touch *)
(* LOC = "X24/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011000011001)
) lut_24_22 (
    .O(x24_y22),
    .I0(x22_y23),
    .I1(x21_y20),
    .I2(x22_y22),
    .I3(x21_y25)
);

(* keep, dont_touch *)
(* LOC = "X25/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000011010010)
) lut_25_22 (
    .O(x25_y22),
    .I0(x23_y27),
    .I1(1'b0),
    .I2(x22_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X26/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110100111110)
) lut_26_22 (
    .O(x26_y22),
    .I0(x23_y24),
    .I1(x24_y22),
    .I2(x24_y17),
    .I3(x23_y18)
);

(* keep, dont_touch *)
(* LOC = "X27/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101001000110)
) lut_27_22 (
    .O(x27_y22),
    .I0(x24_y24),
    .I1(x24_y19),
    .I2(x24_y26),
    .I3(x24_y19)
);

(* keep, dont_touch *)
(* LOC = "X28/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011101111011)
) lut_28_22 (
    .O(x28_y22),
    .I0(x25_y19),
    .I1(x26_y26),
    .I2(x26_y24),
    .I3(x25_y27)
);

(* keep, dont_touch *)
(* LOC = "X29/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101001000010)
) lut_29_22 (
    .O(x29_y22),
    .I0(x27_y18),
    .I1(x26_y21),
    .I2(1'b0),
    .I3(x27_y20)
);

(* keep, dont_touch *)
(* LOC = "X30/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011000110100)
) lut_30_22 (
    .O(x30_y22),
    .I0(x28_y20),
    .I1(x28_y20),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X31/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110101101111)
) lut_31_22 (
    .O(x31_y22),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x29_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X32/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001100100010)
) lut_32_22 (
    .O(x32_y22),
    .I0(x30_y22),
    .I1(1'b0),
    .I2(x30_y24),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X33/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001000000111)
) lut_33_22 (
    .O(x33_y22),
    .I0(1'b0),
    .I1(x30_y19),
    .I2(x31_y18),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X34/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111101010001)
) lut_34_22 (
    .O(x34_y22),
    .I0(x32_y23),
    .I1(x32_y27),
    .I2(1'b0),
    .I3(x32_y21)
);

(* keep, dont_touch *)
(* LOC = "X35/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100000010011)
) lut_35_22 (
    .O(x35_y22),
    .I0(x33_y17),
    .I1(x32_y27),
    .I2(1'b0),
    .I3(x32_y17)
);

(* keep, dont_touch *)
(* LOC = "X36/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110000100110)
) lut_36_22 (
    .O(x36_y22),
    .I0(x33_y24),
    .I1(x34_y27),
    .I2(x34_y26),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X37/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001010011011)
) lut_37_22 (
    .O(x37_y22),
    .I0(x34_y27),
    .I1(x34_y20),
    .I2(x35_y25),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X38/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010100011010)
) lut_38_22 (
    .O(x38_y22),
    .I0(x35_y21),
    .I1(1'b0),
    .I2(x35_y25),
    .I3(x36_y21)
);

(* keep, dont_touch *)
(* LOC = "X39/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101100000010)
) lut_39_22 (
    .O(x39_y22),
    .I0(x36_y25),
    .I1(x36_y23),
    .I2(x36_y25),
    .I3(x37_y24)
);

(* keep, dont_touch *)
(* LOC = "X40/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000101111000)
) lut_40_22 (
    .O(x40_y22),
    .I0(x38_y20),
    .I1(x38_y19),
    .I2(1'b0),
    .I3(x37_y27)
);

(* keep, dont_touch *)
(* LOC = "X41/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011101011111)
) lut_41_22 (
    .O(x41_y22),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x38_y27),
    .I3(x38_y19)
);

(* keep, dont_touch *)
(* LOC = "X42/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110011000100)
) lut_42_22 (
    .O(x42_y22),
    .I0(1'b0),
    .I1(x39_y17),
    .I2(x39_y17),
    .I3(x40_y23)
);

(* keep, dont_touch *)
(* LOC = "X43/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001011100110)
) lut_43_22 (
    .O(x43_y22),
    .I0(x41_y26),
    .I1(1'b0),
    .I2(x41_y27),
    .I3(x40_y20)
);

(* keep, dont_touch *)
(* LOC = "X44/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010111011101)
) lut_44_22 (
    .O(x44_y22),
    .I0(1'b0),
    .I1(x41_y20),
    .I2(1'b0),
    .I3(x42_y20)
);

(* keep, dont_touch *)
(* LOC = "X45/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101101011110)
) lut_45_22 (
    .O(x45_y22),
    .I0(x42_y20),
    .I1(x43_y25),
    .I2(x43_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X46/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101001101000)
) lut_46_22 (
    .O(x46_y22),
    .I0(x44_y25),
    .I1(1'b0),
    .I2(x43_y20),
    .I3(x43_y26)
);

(* keep, dont_touch *)
(* LOC = "X47/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110000000110)
) lut_47_22 (
    .O(x47_y22),
    .I0(x44_y26),
    .I1(x44_y24),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X48/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110000110000)
) lut_48_22 (
    .O(x48_y22),
    .I0(x45_y26),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x46_y24)
);

(* keep, dont_touch *)
(* LOC = "X49/Y22" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010110001011)
) lut_49_22 (
    .O(x49_y22),
    .I0(x47_y24),
    .I1(x46_y22),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X0/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001111001010)
) lut_0_23 (
    .O(x0_y23),
    .I0(1'b0),
    .I1(in7),
    .I2(in3),
    .I3(in4)
);

(* keep, dont_touch *)
(* LOC = "X1/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100011000111)
) lut_1_23 (
    .O(x1_y23),
    .I0(1'b0),
    .I1(in9),
    .I2(in5),
    .I3(in3)
);

(* keep, dont_touch *)
(* LOC = "X2/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110101000101)
) lut_2_23 (
    .O(x2_y23),
    .I0(in0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X3/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011110100011)
) lut_3_23 (
    .O(x3_y23),
    .I0(1'b0),
    .I1(in8),
    .I2(x1_y28),
    .I3(in8)
);

(* keep, dont_touch *)
(* LOC = "X4/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110110011001)
) lut_4_23 (
    .O(x4_y23),
    .I0(x1_y18),
    .I1(x2_y18),
    .I2(x2_y19),
    .I3(x2_y22)
);

(* keep, dont_touch *)
(* LOC = "X5/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000010011101)
) lut_5_23 (
    .O(x5_y23),
    .I0(1'b0),
    .I1(x2_y21),
    .I2(x2_y26),
    .I3(x2_y20)
);

(* keep, dont_touch *)
(* LOC = "X6/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011000011101)
) lut_6_23 (
    .O(x6_y23),
    .I0(x3_y20),
    .I1(x3_y20),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X7/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010111010010)
) lut_7_23 (
    .O(x7_y23),
    .I0(x5_y28),
    .I1(x4_y19),
    .I2(x5_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X8/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000100110111)
) lut_8_23 (
    .O(x8_y23),
    .I0(x5_y20),
    .I1(x6_y20),
    .I2(x6_y20),
    .I3(x5_y20)
);

(* keep, dont_touch *)
(* LOC = "X9/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110001001101)
) lut_9_23 (
    .O(x9_y23),
    .I0(x7_y25),
    .I1(x6_y22),
    .I2(x6_y20),
    .I3(x5_y20)
);

(* keep, dont_touch *)
(* LOC = "X10/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000101110100)
) lut_10_23 (
    .O(x10_y23),
    .I0(x7_y20),
    .I1(x8_y20),
    .I2(x8_y23),
    .I3(x8_y28)
);

(* keep, dont_touch *)
(* LOC = "X11/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100000010101)
) lut_11_23 (
    .O(x11_y23),
    .I0(x8_y19),
    .I1(x9_y27),
    .I2(x9_y27),
    .I3(x8_y20)
);

(* keep, dont_touch *)
(* LOC = "X12/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101001010001)
) lut_12_23 (
    .O(x12_y23),
    .I0(1'b0),
    .I1(x10_y24),
    .I2(x9_y19),
    .I3(x10_y18)
);

(* keep, dont_touch *)
(* LOC = "X13/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001111100101)
) lut_13_23 (
    .O(x13_y23),
    .I0(x11_y21),
    .I1(x10_y19),
    .I2(x10_y26),
    .I3(x11_y20)
);

(* keep, dont_touch *)
(* LOC = "X14/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000001110010)
) lut_14_23 (
    .O(x14_y23),
    .I0(x11_y19),
    .I1(x11_y28),
    .I2(x11_y23),
    .I3(x11_y26)
);

(* keep, dont_touch *)
(* LOC = "X15/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001101001000)
) lut_15_23 (
    .O(x15_y23),
    .I0(x13_y22),
    .I1(x13_y23),
    .I2(1'b0),
    .I3(x12_y24)
);

(* keep, dont_touch *)
(* LOC = "X16/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011001011011)
) lut_16_23 (
    .O(x16_y23),
    .I0(x13_y27),
    .I1(x13_y20),
    .I2(x14_y28),
    .I3(x13_y27)
);

(* keep, dont_touch *)
(* LOC = "X17/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101001101000)
) lut_17_23 (
    .O(x17_y23),
    .I0(x15_y19),
    .I1(x14_y20),
    .I2(1'b0),
    .I3(x15_y27)
);

(* keep, dont_touch *)
(* LOC = "X18/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000011110011)
) lut_18_23 (
    .O(x18_y23),
    .I0(1'b0),
    .I1(x16_y19),
    .I2(x15_y18),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X19/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011110001110)
) lut_19_23 (
    .O(x19_y23),
    .I0(x16_y21),
    .I1(1'b0),
    .I2(x16_y26),
    .I3(x17_y22)
);

(* keep, dont_touch *)
(* LOC = "X20/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101011001111)
) lut_20_23 (
    .O(x20_y23),
    .I0(x17_y21),
    .I1(x17_y22),
    .I2(1'b0),
    .I3(x17_y27)
);

(* keep, dont_touch *)
(* LOC = "X21/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110111101011)
) lut_21_23 (
    .O(x21_y23),
    .I0(x19_y24),
    .I1(x19_y26),
    .I2(x19_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X22/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010001100011)
) lut_22_23 (
    .O(x22_y23),
    .I0(x19_y23),
    .I1(x20_y25),
    .I2(x20_y24),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X23/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100111010101)
) lut_23_23 (
    .O(x23_y23),
    .I0(x20_y22),
    .I1(x21_y22),
    .I2(x21_y19),
    .I3(x21_y24)
);

(* keep, dont_touch *)
(* LOC = "X24/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000011101100)
) lut_24_23 (
    .O(x24_y23),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x22_y22)
);

(* keep, dont_touch *)
(* LOC = "X25/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001001001000)
) lut_25_23 (
    .O(x25_y23),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x22_y23),
    .I3(x23_y20)
);

(* keep, dont_touch *)
(* LOC = "X26/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110111100010)
) lut_26_23 (
    .O(x26_y23),
    .I0(x24_y23),
    .I1(x23_y26),
    .I2(x23_y18),
    .I3(x23_y28)
);

(* keep, dont_touch *)
(* LOC = "X27/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010100001111)
) lut_27_23 (
    .O(x27_y23),
    .I0(1'b0),
    .I1(x25_y19),
    .I2(x24_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X28/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110011011001)
) lut_28_23 (
    .O(x28_y23),
    .I0(x25_y23),
    .I1(x26_y20),
    .I2(x26_y20),
    .I3(x26_y27)
);

(* keep, dont_touch *)
(* LOC = "X29/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101100110010)
) lut_29_23 (
    .O(x29_y23),
    .I0(1'b0),
    .I1(x26_y19),
    .I2(1'b0),
    .I3(x27_y18)
);

(* keep, dont_touch *)
(* LOC = "X30/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111100010110)
) lut_30_23 (
    .O(x30_y23),
    .I0(x28_y18),
    .I1(x28_y20),
    .I2(1'b0),
    .I3(x27_y23)
);

(* keep, dont_touch *)
(* LOC = "X31/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101101011010)
) lut_31_23 (
    .O(x31_y23),
    .I0(x29_y19),
    .I1(1'b0),
    .I2(x29_y25),
    .I3(x28_y19)
);

(* keep, dont_touch *)
(* LOC = "X32/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100101100101)
) lut_32_23 (
    .O(x32_y23),
    .I0(1'b0),
    .I1(x30_y22),
    .I2(x30_y23),
    .I3(x29_y21)
);

(* keep, dont_touch *)
(* LOC = "X33/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101110100100)
) lut_33_23 (
    .O(x33_y23),
    .I0(x31_y23),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x31_y23)
);

(* keep, dont_touch *)
(* LOC = "X34/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110100011100)
) lut_34_23 (
    .O(x34_y23),
    .I0(1'b0),
    .I1(x31_y22),
    .I2(x31_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X35/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001001110000)
) lut_35_23 (
    .O(x35_y23),
    .I0(x32_y21),
    .I1(x32_y27),
    .I2(1'b0),
    .I3(x33_y23)
);

(* keep, dont_touch *)
(* LOC = "X36/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111001110011)
) lut_36_23 (
    .O(x36_y23),
    .I0(1'b0),
    .I1(x34_y19),
    .I2(x33_y24),
    .I3(x34_y26)
);

(* keep, dont_touch *)
(* LOC = "X37/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111111011001)
) lut_37_23 (
    .O(x37_y23),
    .I0(1'b0),
    .I1(x35_y19),
    .I2(x34_y28),
    .I3(x35_y26)
);

(* keep, dont_touch *)
(* LOC = "X38/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010001000001)
) lut_38_23 (
    .O(x38_y23),
    .I0(x35_y23),
    .I1(x36_y19),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X39/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100000000110)
) lut_39_23 (
    .O(x39_y23),
    .I0(1'b0),
    .I1(x37_y22),
    .I2(x37_y24),
    .I3(x36_y23)
);

(* keep, dont_touch *)
(* LOC = "X40/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011101011001)
) lut_40_23 (
    .O(x40_y23),
    .I0(x37_y21),
    .I1(x38_y23),
    .I2(1'b0),
    .I3(x38_y21)
);

(* keep, dont_touch *)
(* LOC = "X41/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111110001110)
) lut_41_23 (
    .O(x41_y23),
    .I0(x39_y27),
    .I1(x39_y24),
    .I2(x39_y25),
    .I3(x38_y28)
);

(* keep, dont_touch *)
(* LOC = "X42/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000100000000)
) lut_42_23 (
    .O(x42_y23),
    .I0(x39_y18),
    .I1(x40_y18),
    .I2(x40_y22),
    .I3(x40_y22)
);

(* keep, dont_touch *)
(* LOC = "X43/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000001001010)
) lut_43_23 (
    .O(x43_y23),
    .I0(x40_y25),
    .I1(x40_y22),
    .I2(x41_y19),
    .I3(x40_y26)
);

(* keep, dont_touch *)
(* LOC = "X44/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011110011101)
) lut_44_23 (
    .O(x44_y23),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x42_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X45/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100001000101)
) lut_45_23 (
    .O(x45_y23),
    .I0(x43_y23),
    .I1(x43_y27),
    .I2(x42_y19),
    .I3(x43_y20)
);

(* keep, dont_touch *)
(* LOC = "X46/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000010000101)
) lut_46_23 (
    .O(x46_y23),
    .I0(x44_y20),
    .I1(1'b0),
    .I2(x44_y18),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X47/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100000011000)
) lut_47_23 (
    .O(x47_y23),
    .I0(x44_y27),
    .I1(1'b0),
    .I2(x44_y18),
    .I3(x44_y28)
);

(* keep, dont_touch *)
(* LOC = "X48/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010110010100)
) lut_48_23 (
    .O(x48_y23),
    .I0(x45_y28),
    .I1(x46_y19),
    .I2(1'b0),
    .I3(x46_y26)
);

(* keep, dont_touch *)
(* LOC = "X49/Y23" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000011110110)
) lut_49_23 (
    .O(x49_y23),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x47_y24),
    .I3(x47_y23)
);

(* keep, dont_touch *)
(* LOC = "X0/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011010110101)
) lut_0_24 (
    .O(x0_y24),
    .I0(in7),
    .I1(1'b0),
    .I2(in1),
    .I3(in3)
);

(* keep, dont_touch *)
(* LOC = "X1/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111100011000)
) lut_1_24 (
    .O(x1_y24),
    .I0(in5),
    .I1(in3),
    .I2(in0),
    .I3(in0)
);

(* keep, dont_touch *)
(* LOC = "X2/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111110110010)
) lut_2_24 (
    .O(x2_y24),
    .I0(in4),
    .I1(in1),
    .I2(in9),
    .I3(in5)
);

(* keep, dont_touch *)
(* LOC = "X3/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111110111001)
) lut_3_24 (
    .O(x3_y24),
    .I0(x1_y23),
    .I1(1'b0),
    .I2(in3),
    .I3(in7)
);

(* keep, dont_touch *)
(* LOC = "X4/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001010011010)
) lut_4_24 (
    .O(x4_y24),
    .I0(x1_y19),
    .I1(x2_y21),
    .I2(1'b0),
    .I3(x2_y21)
);

(* keep, dont_touch *)
(* LOC = "X5/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110000001000)
) lut_5_24 (
    .O(x5_y24),
    .I0(x2_y29),
    .I1(x2_y19),
    .I2(1'b0),
    .I3(x2_y22)
);

(* keep, dont_touch *)
(* LOC = "X6/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100111100111)
) lut_6_24 (
    .O(x6_y24),
    .I0(x3_y21),
    .I1(x4_y21),
    .I2(x3_y20),
    .I3(x4_y26)
);

(* keep, dont_touch *)
(* LOC = "X7/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100011101001)
) lut_7_24 (
    .O(x7_y24),
    .I0(x5_y19),
    .I1(x4_y19),
    .I2(x5_y24),
    .I3(x5_y20)
);

(* keep, dont_touch *)
(* LOC = "X8/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000100110000)
) lut_8_24 (
    .O(x8_y24),
    .I0(x6_y28),
    .I1(x6_y23),
    .I2(1'b0),
    .I3(x6_y21)
);

(* keep, dont_touch *)
(* LOC = "X9/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000101110011)
) lut_9_24 (
    .O(x9_y24),
    .I0(x6_y19),
    .I1(x6_y22),
    .I2(1'b0),
    .I3(x6_y21)
);

(* keep, dont_touch *)
(* LOC = "X10/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101000011011)
) lut_10_24 (
    .O(x10_y24),
    .I0(1'b0),
    .I1(x7_y21),
    .I2(1'b0),
    .I3(x8_y19)
);

(* keep, dont_touch *)
(* LOC = "X11/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101010100111)
) lut_11_24 (
    .O(x11_y24),
    .I0(x8_y24),
    .I1(1'b0),
    .I2(x8_y26),
    .I3(x9_y25)
);

(* keep, dont_touch *)
(* LOC = "X12/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011111110101)
) lut_12_24 (
    .O(x12_y24),
    .I0(x10_y27),
    .I1(x10_y22),
    .I2(x9_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X13/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101010110100)
) lut_13_24 (
    .O(x13_y24),
    .I0(x11_y19),
    .I1(x10_y19),
    .I2(x10_y21),
    .I3(x11_y22)
);

(* keep, dont_touch *)
(* LOC = "X14/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100010100000)
) lut_14_24 (
    .O(x14_y24),
    .I0(x12_y28),
    .I1(x11_y24),
    .I2(x11_y22),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X15/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101100010111)
) lut_15_24 (
    .O(x15_y24),
    .I0(x12_y26),
    .I1(x12_y23),
    .I2(x12_y19),
    .I3(x13_y19)
);

(* keep, dont_touch *)
(* LOC = "X16/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000011001101)
) lut_16_24 (
    .O(x16_y24),
    .I0(x13_y28),
    .I1(1'b0),
    .I2(x13_y22),
    .I3(x13_y22)
);

(* keep, dont_touch *)
(* LOC = "X17/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110101010101)
) lut_17_24 (
    .O(x17_y24),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X18/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101001011011)
) lut_18_24 (
    .O(x18_y24),
    .I0(x16_y24),
    .I1(x15_y20),
    .I2(x16_y28),
    .I3(x15_y19)
);

(* keep, dont_touch *)
(* LOC = "X19/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111000101111)
) lut_19_24 (
    .O(x19_y24),
    .I0(x17_y27),
    .I1(x16_y20),
    .I2(x17_y25),
    .I3(x16_y20)
);

(* keep, dont_touch *)
(* LOC = "X20/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101001011001)
) lut_20_24 (
    .O(x20_y24),
    .I0(x18_y19),
    .I1(x18_y27),
    .I2(1'b0),
    .I3(x18_y19)
);

(* keep, dont_touch *)
(* LOC = "X21/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111010110111)
) lut_21_24 (
    .O(x21_y24),
    .I0(x18_y24),
    .I1(x18_y28),
    .I2(x19_y21),
    .I3(x18_y23)
);

(* keep, dont_touch *)
(* LOC = "X22/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001010101000)
) lut_22_24 (
    .O(x22_y24),
    .I0(x20_y28),
    .I1(x19_y25),
    .I2(x19_y20),
    .I3(x20_y27)
);

(* keep, dont_touch *)
(* LOC = "X23/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011100110011)
) lut_23_24 (
    .O(x23_y24),
    .I0(x20_y21),
    .I1(x21_y19),
    .I2(x20_y26),
    .I3(x20_y23)
);

(* keep, dont_touch *)
(* LOC = "X24/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101111110011)
) lut_24_24 (
    .O(x24_y24),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x21_y20),
    .I3(x22_y20)
);

(* keep, dont_touch *)
(* LOC = "X25/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001101110111)
) lut_25_24 (
    .O(x25_y24),
    .I0(x22_y29),
    .I1(x22_y28),
    .I2(x22_y26),
    .I3(x23_y22)
);

(* keep, dont_touch *)
(* LOC = "X26/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101100111111)
) lut_26_24 (
    .O(x26_y24),
    .I0(x23_y28),
    .I1(x24_y22),
    .I2(x23_y19),
    .I3(x24_y20)
);

(* keep, dont_touch *)
(* LOC = "X27/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000000011100)
) lut_27_24 (
    .O(x27_y24),
    .I0(x24_y29),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X28/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111001010111)
) lut_28_24 (
    .O(x28_y24),
    .I0(x25_y21),
    .I1(x26_y28),
    .I2(1'b0),
    .I3(x26_y27)
);

(* keep, dont_touch *)
(* LOC = "X29/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011110000100)
) lut_29_24 (
    .O(x29_y24),
    .I0(x27_y26),
    .I1(1'b0),
    .I2(x26_y20),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X30/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001101101100)
) lut_30_24 (
    .O(x30_y24),
    .I0(x28_y25),
    .I1(x28_y22),
    .I2(1'b0),
    .I3(x27_y26)
);

(* keep, dont_touch *)
(* LOC = "X31/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100101101011)
) lut_31_24 (
    .O(x31_y24),
    .I0(x28_y25),
    .I1(x28_y24),
    .I2(x28_y22),
    .I3(x28_y26)
);

(* keep, dont_touch *)
(* LOC = "X32/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000100101100)
) lut_32_24 (
    .O(x32_y24),
    .I0(x29_y20),
    .I1(x29_y19),
    .I2(x29_y23),
    .I3(x30_y20)
);

(* keep, dont_touch *)
(* LOC = "X33/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100000100111)
) lut_33_24 (
    .O(x33_y24),
    .I0(1'b0),
    .I1(x30_y27),
    .I2(x30_y21),
    .I3(x31_y23)
);

(* keep, dont_touch *)
(* LOC = "X34/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101011101100)
) lut_34_24 (
    .O(x34_y24),
    .I0(x32_y26),
    .I1(x31_y26),
    .I2(x31_y24),
    .I3(x31_y27)
);

(* keep, dont_touch *)
(* LOC = "X35/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111100110010)
) lut_35_24 (
    .O(x35_y24),
    .I0(x33_y26),
    .I1(1'b0),
    .I2(x33_y24),
    .I3(x33_y29)
);

(* keep, dont_touch *)
(* LOC = "X36/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010100000101)
) lut_36_24 (
    .O(x36_y24),
    .I0(x33_y28),
    .I1(x34_y19),
    .I2(x34_y19),
    .I3(x33_y28)
);

(* keep, dont_touch *)
(* LOC = "X37/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011000000110)
) lut_37_24 (
    .O(x37_y24),
    .I0(x35_y27),
    .I1(x35_y24),
    .I2(x34_y23),
    .I3(x34_y19)
);

(* keep, dont_touch *)
(* LOC = "X38/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100001010001)
) lut_38_24 (
    .O(x38_y24),
    .I0(x35_y27),
    .I1(x35_y27),
    .I2(x36_y20),
    .I3(x35_y19)
);

(* keep, dont_touch *)
(* LOC = "X39/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101100100111)
) lut_39_24 (
    .O(x39_y24),
    .I0(x36_y24),
    .I1(x37_y24),
    .I2(x37_y26),
    .I3(x37_y27)
);

(* keep, dont_touch *)
(* LOC = "X40/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111001011000)
) lut_40_24 (
    .O(x40_y24),
    .I0(x38_y29),
    .I1(x37_y22),
    .I2(x37_y22),
    .I3(x37_y25)
);

(* keep, dont_touch *)
(* LOC = "X41/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000110000111)
) lut_41_24 (
    .O(x41_y24),
    .I0(x39_y24),
    .I1(1'b0),
    .I2(x38_y27),
    .I3(x39_y24)
);

(* keep, dont_touch *)
(* LOC = "X42/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000110111110)
) lut_42_24 (
    .O(x42_y24),
    .I0(1'b0),
    .I1(x39_y25),
    .I2(1'b0),
    .I3(x40_y25)
);

(* keep, dont_touch *)
(* LOC = "X43/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110000101111)
) lut_43_24 (
    .O(x43_y24),
    .I0(x41_y29),
    .I1(x40_y22),
    .I2(x40_y19),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X44/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000101111111)
) lut_44_24 (
    .O(x44_y24),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x42_y23),
    .I3(x41_y23)
);

(* keep, dont_touch *)
(* LOC = "X45/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010101111101)
) lut_45_24 (
    .O(x45_y24),
    .I0(1'b0),
    .I1(x43_y28),
    .I2(x43_y26),
    .I3(x43_y29)
);

(* keep, dont_touch *)
(* LOC = "X46/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100001000010)
) lut_46_24 (
    .O(x46_y24),
    .I0(x43_y23),
    .I1(x43_y19),
    .I2(1'b0),
    .I3(x43_y28)
);

(* keep, dont_touch *)
(* LOC = "X47/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111011010001)
) lut_47_24 (
    .O(x47_y24),
    .I0(x45_y25),
    .I1(x45_y25),
    .I2(x44_y20),
    .I3(x45_y29)
);

(* keep, dont_touch *)
(* LOC = "X48/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101001010101)
) lut_48_24 (
    .O(x48_y24),
    .I0(x46_y21),
    .I1(x46_y20),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X49/Y24" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000000111010)
) lut_49_24 (
    .O(x49_y24),
    .I0(x47_y24),
    .I1(x46_y23),
    .I2(x46_y24),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X0/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011101111110)
) lut_0_25 (
    .O(x0_y25),
    .I0(in9),
    .I1(in0),
    .I2(in9),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X1/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101001110110)
) lut_1_25 (
    .O(x1_y25),
    .I0(in8),
    .I1(in5),
    .I2(in4),
    .I3(in7)
);

(* keep, dont_touch *)
(* LOC = "X2/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100100100110)
) lut_2_25 (
    .O(x2_y25),
    .I0(in5),
    .I1(in4),
    .I2(in5),
    .I3(in0)
);

(* keep, dont_touch *)
(* LOC = "X3/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001010011111)
) lut_3_25 (
    .O(x3_y25),
    .I0(x1_y29),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X4/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110111100011)
) lut_4_25 (
    .O(x4_y25),
    .I0(x2_y28),
    .I1(x1_y29),
    .I2(1'b0),
    .I3(x1_y25)
);

(* keep, dont_touch *)
(* LOC = "X5/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100101010110)
) lut_5_25 (
    .O(x5_y25),
    .I0(1'b0),
    .I1(x3_y23),
    .I2(1'b0),
    .I3(x2_y29)
);

(* keep, dont_touch *)
(* LOC = "X6/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101101110010)
) lut_6_25 (
    .O(x6_y25),
    .I0(x3_y30),
    .I1(x3_y24),
    .I2(x3_y20),
    .I3(x4_y25)
);

(* keep, dont_touch *)
(* LOC = "X7/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101101010110)
) lut_7_25 (
    .O(x7_y25),
    .I0(1'b0),
    .I1(x5_y26),
    .I2(1'b0),
    .I3(x5_y25)
);

(* keep, dont_touch *)
(* LOC = "X8/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100001010111)
) lut_8_25 (
    .O(x8_y25),
    .I0(x5_y21),
    .I1(1'b0),
    .I2(x5_y29),
    .I3(x5_y29)
);

(* keep, dont_touch *)
(* LOC = "X9/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100101100000)
) lut_9_25 (
    .O(x9_y25),
    .I0(x6_y30),
    .I1(1'b0),
    .I2(x5_y29),
    .I3(x5_y29)
);

(* keep, dont_touch *)
(* LOC = "X10/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001011100010)
) lut_10_25 (
    .O(x10_y25),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x8_y26)
);

(* keep, dont_touch *)
(* LOC = "X11/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101111010111)
) lut_11_25 (
    .O(x11_y25),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x8_y28)
);

(* keep, dont_touch *)
(* LOC = "X12/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010000000101)
) lut_12_25 (
    .O(x12_y25),
    .I0(x10_y29),
    .I1(x10_y29),
    .I2(x10_y20),
    .I3(x9_y26)
);

(* keep, dont_touch *)
(* LOC = "X13/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011111111011)
) lut_13_25 (
    .O(x13_y25),
    .I0(1'b0),
    .I1(x11_y28),
    .I2(x10_y25),
    .I3(x11_y26)
);

(* keep, dont_touch *)
(* LOC = "X14/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001101000001)
) lut_14_25 (
    .O(x14_y25),
    .I0(1'b0),
    .I1(x12_y24),
    .I2(1'b0),
    .I3(x11_y26)
);

(* keep, dont_touch *)
(* LOC = "X15/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011111110110)
) lut_15_25 (
    .O(x15_y25),
    .I0(x12_y26),
    .I1(x12_y21),
    .I2(x13_y21),
    .I3(x13_y30)
);

(* keep, dont_touch *)
(* LOC = "X16/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010001001110)
) lut_16_25 (
    .O(x16_y25),
    .I0(x13_y28),
    .I1(1'b0),
    .I2(x14_y26),
    .I3(x13_y29)
);

(* keep, dont_touch *)
(* LOC = "X17/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000010100010)
) lut_17_25 (
    .O(x17_y25),
    .I0(x15_y23),
    .I1(x15_y27),
    .I2(x15_y29),
    .I3(x15_y29)
);

(* keep, dont_touch *)
(* LOC = "X18/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111010100110)
) lut_18_25 (
    .O(x18_y25),
    .I0(x15_y30),
    .I1(1'b0),
    .I2(x16_y30),
    .I3(x15_y25)
);

(* keep, dont_touch *)
(* LOC = "X19/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100000111011)
) lut_19_25 (
    .O(x19_y25),
    .I0(1'b0),
    .I1(x17_y29),
    .I2(x17_y27),
    .I3(x16_y20)
);

(* keep, dont_touch *)
(* LOC = "X20/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000101101000)
) lut_20_25 (
    .O(x20_y25),
    .I0(x18_y23),
    .I1(x17_y28),
    .I2(x18_y21),
    .I3(x18_y22)
);

(* keep, dont_touch *)
(* LOC = "X21/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101101001110)
) lut_21_25 (
    .O(x21_y25),
    .I0(x18_y26),
    .I1(x18_y27),
    .I2(x19_y28),
    .I3(x19_y29)
);

(* keep, dont_touch *)
(* LOC = "X22/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001000011101)
) lut_22_25 (
    .O(x22_y25),
    .I0(x20_y23),
    .I1(x19_y28),
    .I2(x20_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X23/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110001000010)
) lut_23_25 (
    .O(x23_y25),
    .I0(x20_y22),
    .I1(x21_y25),
    .I2(1'b0),
    .I3(x20_y25)
);

(* keep, dont_touch *)
(* LOC = "X24/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000001100011)
) lut_24_25 (
    .O(x24_y25),
    .I0(x21_y24),
    .I1(x22_y26),
    .I2(1'b0),
    .I3(x22_y28)
);

(* keep, dont_touch *)
(* LOC = "X25/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110001001111)
) lut_25_25 (
    .O(x25_y25),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x23_y22),
    .I3(x23_y24)
);

(* keep, dont_touch *)
(* LOC = "X26/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100000001110)
) lut_26_25 (
    .O(x26_y25),
    .I0(x23_y22),
    .I1(x24_y20),
    .I2(x23_y22),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X27/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001010110010)
) lut_27_25 (
    .O(x27_y25),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x25_y20)
);

(* keep, dont_touch *)
(* LOC = "X28/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010110010100)
) lut_28_25 (
    .O(x28_y25),
    .I0(x26_y24),
    .I1(x25_y28),
    .I2(x25_y28),
    .I3(x26_y24)
);

(* keep, dont_touch *)
(* LOC = "X29/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000011101011)
) lut_29_25 (
    .O(x29_y25),
    .I0(x26_y23),
    .I1(x27_y20),
    .I2(x26_y25),
    .I3(x26_y29)
);

(* keep, dont_touch *)
(* LOC = "X30/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100110111010)
) lut_30_25 (
    .O(x30_y25),
    .I0(x27_y26),
    .I1(x27_y26),
    .I2(x28_y23),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X31/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000110101000)
) lut_31_25 (
    .O(x31_y25),
    .I0(x29_y28),
    .I1(1'b0),
    .I2(x29_y22),
    .I3(x28_y29)
);

(* keep, dont_touch *)
(* LOC = "X32/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111011011100)
) lut_32_25 (
    .O(x32_y25),
    .I0(x30_y28),
    .I1(1'b0),
    .I2(x30_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X33/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111111101011)
) lut_33_25 (
    .O(x33_y25),
    .I0(x30_y23),
    .I1(x31_y23),
    .I2(x31_y29),
    .I3(x30_y23)
);

(* keep, dont_touch *)
(* LOC = "X34/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001011111110)
) lut_34_25 (
    .O(x34_y25),
    .I0(x32_y25),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x31_y25)
);

(* keep, dont_touch *)
(* LOC = "X35/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001011011000)
) lut_35_25 (
    .O(x35_y25),
    .I0(1'b0),
    .I1(x32_y29),
    .I2(x33_y21),
    .I3(x33_y24)
);

(* keep, dont_touch *)
(* LOC = "X36/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110100001010)
) lut_36_25 (
    .O(x36_y25),
    .I0(1'b0),
    .I1(x34_y29),
    .I2(x33_y26),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X37/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110011001011)
) lut_37_25 (
    .O(x37_y25),
    .I0(x35_y29),
    .I1(x34_y30),
    .I2(x35_y28),
    .I3(x34_y26)
);

(* keep, dont_touch *)
(* LOC = "X38/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110000001010)
) lut_38_25 (
    .O(x38_y25),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x35_y22),
    .I3(x36_y20)
);

(* keep, dont_touch *)
(* LOC = "X39/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100010111111)
) lut_39_25 (
    .O(x39_y25),
    .I0(x36_y25),
    .I1(x36_y22),
    .I2(x36_y28),
    .I3(x37_y27)
);

(* keep, dont_touch *)
(* LOC = "X40/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010101011100)
) lut_40_25 (
    .O(x40_y25),
    .I0(x38_y30),
    .I1(1'b0),
    .I2(x38_y27),
    .I3(x37_y23)
);

(* keep, dont_touch *)
(* LOC = "X41/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100010101011)
) lut_41_25 (
    .O(x41_y25),
    .I0(x39_y25),
    .I1(x38_y20),
    .I2(1'b0),
    .I3(x39_y23)
);

(* keep, dont_touch *)
(* LOC = "X42/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101110001101)
) lut_42_25 (
    .O(x42_y25),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x39_y29),
    .I3(x40_y25)
);

(* keep, dont_touch *)
(* LOC = "X43/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110000011001)
) lut_43_25 (
    .O(x43_y25),
    .I0(x41_y23),
    .I1(x40_y30),
    .I2(1'b0),
    .I3(x41_y25)
);

(* keep, dont_touch *)
(* LOC = "X44/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110100010111)
) lut_44_25 (
    .O(x44_y25),
    .I0(x41_y21),
    .I1(x41_y23),
    .I2(x41_y23),
    .I3(x42_y23)
);

(* keep, dont_touch *)
(* LOC = "X45/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001011011111)
) lut_45_25 (
    .O(x45_y25),
    .I0(x43_y28),
    .I1(x43_y28),
    .I2(x43_y29),
    .I3(x43_y22)
);

(* keep, dont_touch *)
(* LOC = "X46/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100000111000)
) lut_46_25 (
    .O(x46_y25),
    .I0(x44_y23),
    .I1(x43_y29),
    .I2(x44_y30),
    .I3(x43_y27)
);

(* keep, dont_touch *)
(* LOC = "X47/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110010111011)
) lut_47_25 (
    .O(x47_y25),
    .I0(1'b0),
    .I1(x44_y25),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X48/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100101011101)
) lut_48_25 (
    .O(x48_y25),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x45_y24),
    .I3(x46_y21)
);

(* keep, dont_touch *)
(* LOC = "X49/Y25" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100001111100)
) lut_49_25 (
    .O(x49_y25),
    .I0(x47_y23),
    .I1(1'b0),
    .I2(x46_y29),
    .I3(x47_y26)
);

(* keep, dont_touch *)
(* LOC = "X0/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101000000111)
) lut_0_26 (
    .O(x0_y26),
    .I0(in9),
    .I1(1'b0),
    .I2(1'b0),
    .I3(in1)
);

(* keep, dont_touch *)
(* LOC = "X1/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001001000100)
) lut_1_26 (
    .O(x1_y26),
    .I0(1'b0),
    .I1(in1),
    .I2(in8),
    .I3(in3)
);

(* keep, dont_touch *)
(* LOC = "X2/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000010001010)
) lut_2_26 (
    .O(x2_y26),
    .I0(in2),
    .I1(1'b0),
    .I2(in8),
    .I3(in3)
);

(* keep, dont_touch *)
(* LOC = "X3/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101010011101)
) lut_3_26 (
    .O(x3_y26),
    .I0(in0),
    .I1(1'b0),
    .I2(x1_y26),
    .I3(in8)
);

(* keep, dont_touch *)
(* LOC = "X4/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101100110001)
) lut_4_26 (
    .O(x4_y26),
    .I0(1'b0),
    .I1(x2_y28),
    .I2(1'b0),
    .I3(x2_y27)
);

(* keep, dont_touch *)
(* LOC = "X5/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111011011000)
) lut_5_26 (
    .O(x5_y26),
    .I0(1'b0),
    .I1(x3_y28),
    .I2(x3_y27),
    .I3(x3_y31)
);

(* keep, dont_touch *)
(* LOC = "X6/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110001001100)
) lut_6_26 (
    .O(x6_y26),
    .I0(1'b0),
    .I1(x3_y21),
    .I2(x4_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X7/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000000000011)
) lut_7_26 (
    .O(x7_y26),
    .I0(x5_y30),
    .I1(x4_y29),
    .I2(x4_y30),
    .I3(x5_y31)
);

(* keep, dont_touch *)
(* LOC = "X8/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010001010011)
) lut_8_26 (
    .O(x8_y26),
    .I0(x6_y30),
    .I1(x6_y22),
    .I2(x6_y29),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X9/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010100000100)
) lut_9_26 (
    .O(x9_y26),
    .I0(x7_y23),
    .I1(x7_y28),
    .I2(x6_y29),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X10/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001101100010)
) lut_10_26 (
    .O(x10_y26),
    .I0(x8_y22),
    .I1(x8_y29),
    .I2(x8_y28),
    .I3(x8_y23)
);

(* keep, dont_touch *)
(* LOC = "X11/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101011010011)
) lut_11_26 (
    .O(x11_y26),
    .I0(x8_y26),
    .I1(x9_y31),
    .I2(x9_y28),
    .I3(x9_y29)
);

(* keep, dont_touch *)
(* LOC = "X12/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011011101111)
) lut_12_26 (
    .O(x12_y26),
    .I0(x9_y23),
    .I1(x10_y31),
    .I2(1'b0),
    .I3(x9_y28)
);

(* keep, dont_touch *)
(* LOC = "X13/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011010001011)
) lut_13_26 (
    .O(x13_y26),
    .I0(x11_y30),
    .I1(x10_y24),
    .I2(x10_y23),
    .I3(x10_y30)
);

(* keep, dont_touch *)
(* LOC = "X14/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001010010101)
) lut_14_26 (
    .O(x14_y26),
    .I0(x12_y23),
    .I1(x12_y21),
    .I2(x11_y25),
    .I3(x11_y25)
);

(* keep, dont_touch *)
(* LOC = "X15/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100010100011)
) lut_15_26 (
    .O(x15_y26),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x13_y31)
);

(* keep, dont_touch *)
(* LOC = "X16/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100001000100)
) lut_16_26 (
    .O(x16_y26),
    .I0(x14_y25),
    .I1(x14_y21),
    .I2(x13_y21),
    .I3(x13_y28)
);

(* keep, dont_touch *)
(* LOC = "X17/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000010010001)
) lut_17_26 (
    .O(x17_y26),
    .I0(x14_y31),
    .I1(x15_y30),
    .I2(x14_y25),
    .I3(x14_y26)
);

(* keep, dont_touch *)
(* LOC = "X18/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001000110101)
) lut_18_26 (
    .O(x18_y26),
    .I0(1'b0),
    .I1(x16_y26),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X19/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110011001101)
) lut_19_26 (
    .O(x19_y26),
    .I0(1'b0),
    .I1(x17_y21),
    .I2(1'b0),
    .I3(x17_y31)
);

(* keep, dont_touch *)
(* LOC = "X20/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000011101010)
) lut_20_26 (
    .O(x20_y26),
    .I0(x17_y27),
    .I1(x17_y23),
    .I2(x18_y30),
    .I3(x17_y22)
);

(* keep, dont_touch *)
(* LOC = "X21/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010101110100)
) lut_21_26 (
    .O(x21_y26),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x19_y21),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X22/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100110100110)
) lut_22_26 (
    .O(x22_y26),
    .I0(x19_y22),
    .I1(1'b0),
    .I2(x20_y29),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X23/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110011100111)
) lut_23_26 (
    .O(x23_y26),
    .I0(x20_y27),
    .I1(x20_y28),
    .I2(x20_y27),
    .I3(x21_y26)
);

(* keep, dont_touch *)
(* LOC = "X24/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000101110000)
) lut_24_26 (
    .O(x24_y26),
    .I0(1'b0),
    .I1(x22_y22),
    .I2(1'b0),
    .I3(x22_y31)
);

(* keep, dont_touch *)
(* LOC = "X25/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111101000010)
) lut_25_26 (
    .O(x25_y26),
    .I0(x22_y30),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x23_y30)
);

(* keep, dont_touch *)
(* LOC = "X26/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000110111111)
) lut_26_26 (
    .O(x26_y26),
    .I0(1'b0),
    .I1(x23_y27),
    .I2(x24_y21),
    .I3(x23_y25)
);

(* keep, dont_touch *)
(* LOC = "X27/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100000111111)
) lut_27_26 (
    .O(x27_y26),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x24_y22),
    .I3(x24_y25)
);

(* keep, dont_touch *)
(* LOC = "X28/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001001000001)
) lut_28_26 (
    .O(x28_y26),
    .I0(x25_y23),
    .I1(x25_y27),
    .I2(x26_y31),
    .I3(x25_y27)
);

(* keep, dont_touch *)
(* LOC = "X29/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001111111001)
) lut_29_26 (
    .O(x29_y26),
    .I0(x26_y29),
    .I1(x27_y21),
    .I2(1'b0),
    .I3(x27_y24)
);

(* keep, dont_touch *)
(* LOC = "X30/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110101000000)
) lut_30_26 (
    .O(x30_y26),
    .I0(x28_y29),
    .I1(x28_y30),
    .I2(x27_y25),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X31/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000011001100)
) lut_31_26 (
    .O(x31_y26),
    .I0(x28_y24),
    .I1(x28_y30),
    .I2(x29_y25),
    .I3(x29_y22)
);

(* keep, dont_touch *)
(* LOC = "X32/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000110010111)
) lut_32_26 (
    .O(x32_y26),
    .I0(x30_y28),
    .I1(x30_y30),
    .I2(x29_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X33/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000010110010)
) lut_33_26 (
    .O(x33_y26),
    .I0(1'b0),
    .I1(x30_y22),
    .I2(x31_y22),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X34/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011111110101)
) lut_34_26 (
    .O(x34_y26),
    .I0(x32_y30),
    .I1(x32_y23),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X35/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100111111111)
) lut_35_26 (
    .O(x35_y26),
    .I0(x33_y22),
    .I1(x32_y28),
    .I2(x32_y26),
    .I3(x33_y23)
);

(* keep, dont_touch *)
(* LOC = "X36/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111001010001)
) lut_36_26 (
    .O(x36_y26),
    .I0(x33_y27),
    .I1(x33_y27),
    .I2(x33_y22),
    .I3(x34_y26)
);

(* keep, dont_touch *)
(* LOC = "X37/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000100001001)
) lut_37_26 (
    .O(x37_y26),
    .I0(x35_y23),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x34_y29)
);

(* keep, dont_touch *)
(* LOC = "X38/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100001010010)
) lut_38_26 (
    .O(x38_y26),
    .I0(1'b0),
    .I1(x35_y24),
    .I2(x35_y30),
    .I3(x35_y27)
);

(* keep, dont_touch *)
(* LOC = "X39/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011001101001)
) lut_39_26 (
    .O(x39_y26),
    .I0(x36_y27),
    .I1(1'b0),
    .I2(x36_y24),
    .I3(x36_y27)
);

(* keep, dont_touch *)
(* LOC = "X40/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011000110100)
) lut_40_26 (
    .O(x40_y26),
    .I0(1'b0),
    .I1(x38_y24),
    .I2(1'b0),
    .I3(x37_y21)
);

(* keep, dont_touch *)
(* LOC = "X41/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000011001001)
) lut_41_26 (
    .O(x41_y26),
    .I0(1'b0),
    .I1(x38_y24),
    .I2(x38_y31),
    .I3(x38_y25)
);

(* keep, dont_touch *)
(* LOC = "X42/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111101100010)
) lut_42_26 (
    .O(x42_y26),
    .I0(x40_y23),
    .I1(x40_y23),
    .I2(x40_y25),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X43/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111110011101)
) lut_43_26 (
    .O(x43_y26),
    .I0(x41_y28),
    .I1(x40_y30),
    .I2(x40_y26),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X44/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111101010100)
) lut_44_26 (
    .O(x44_y26),
    .I0(x41_y29),
    .I1(x41_y25),
    .I2(x42_y31),
    .I3(x41_y23)
);

(* keep, dont_touch *)
(* LOC = "X45/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010111010010)
) lut_45_26 (
    .O(x45_y26),
    .I0(1'b0),
    .I1(x42_y26),
    .I2(x43_y27),
    .I3(x42_y21)
);

(* keep, dont_touch *)
(* LOC = "X46/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001011111110)
) lut_46_26 (
    .O(x46_y26),
    .I0(x44_y29),
    .I1(x43_y22),
    .I2(x43_y31),
    .I3(x44_y30)
);

(* keep, dont_touch *)
(* LOC = "X47/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100110011111)
) lut_47_26 (
    .O(x47_y26),
    .I0(x44_y28),
    .I1(x45_y26),
    .I2(x44_y27),
    .I3(x44_y23)
);

(* keep, dont_touch *)
(* LOC = "X48/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111011000110)
) lut_48_26 (
    .O(x48_y26),
    .I0(x46_y31),
    .I1(x46_y22),
    .I2(1'b0),
    .I3(x46_y28)
);

(* keep, dont_touch *)
(* LOC = "X49/Y26" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000001110101)
) lut_49_26 (
    .O(x49_y26),
    .I0(x47_y28),
    .I1(x47_y25),
    .I2(x46_y26),
    .I3(x46_y24)
);

(* keep, dont_touch *)
(* LOC = "X0/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001010110100)
) lut_0_27 (
    .O(x0_y27),
    .I0(1'b0),
    .I1(in2),
    .I2(in7),
    .I3(in7)
);

(* keep, dont_touch *)
(* LOC = "X1/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101100010000)
) lut_1_27 (
    .O(x1_y27),
    .I0(1'b0),
    .I1(in7),
    .I2(in7),
    .I3(in4)
);

(* keep, dont_touch *)
(* LOC = "X2/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101011110100)
) lut_2_27 (
    .O(x2_y27),
    .I0(in2),
    .I1(in6),
    .I2(in6),
    .I3(in0)
);

(* keep, dont_touch *)
(* LOC = "X3/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010110011000)
) lut_3_27 (
    .O(x3_y27),
    .I0(x1_y26),
    .I1(in2),
    .I2(in1),
    .I3(in1)
);

(* keep, dont_touch *)
(* LOC = "X4/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101101100000)
) lut_4_27 (
    .O(x4_y27),
    .I0(x1_y31),
    .I1(x1_y22),
    .I2(x1_y27),
    .I3(x2_y23)
);

(* keep, dont_touch *)
(* LOC = "X5/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100100010111)
) lut_5_27 (
    .O(x5_y27),
    .I0(x3_y32),
    .I1(x3_y24),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X6/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100001111111)
) lut_6_27 (
    .O(x6_y27),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x3_y27),
    .I3(x3_y22)
);

(* keep, dont_touch *)
(* LOC = "X7/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100111000110)
) lut_7_27 (
    .O(x7_y27),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x5_y23)
);

(* keep, dont_touch *)
(* LOC = "X8/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101101000111)
) lut_8_27 (
    .O(x8_y27),
    .I0(x6_y22),
    .I1(x6_y30),
    .I2(x6_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X9/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111110010000)
) lut_9_27 (
    .O(x9_y27),
    .I0(x6_y32),
    .I1(x7_y31),
    .I2(x6_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X10/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000110000111)
) lut_10_27 (
    .O(x10_y27),
    .I0(x8_y22),
    .I1(x7_y32),
    .I2(x8_y24),
    .I3(x7_y29)
);

(* keep, dont_touch *)
(* LOC = "X11/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010001011100)
) lut_11_27 (
    .O(x11_y27),
    .I0(x8_y29),
    .I1(x8_y24),
    .I2(x8_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X12/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101011100100)
) lut_12_27 (
    .O(x12_y27),
    .I0(x10_y27),
    .I1(1'b0),
    .I2(x9_y32),
    .I3(x9_y31)
);

(* keep, dont_touch *)
(* LOC = "X13/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110110010100)
) lut_13_27 (
    .O(x13_y27),
    .I0(1'b0),
    .I1(x11_y31),
    .I2(x10_y26),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X14/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101100101111)
) lut_14_27 (
    .O(x14_y27),
    .I0(x12_y28),
    .I1(x12_y31),
    .I2(x12_y31),
    .I3(x11_y22)
);

(* keep, dont_touch *)
(* LOC = "X15/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100011111100)
) lut_15_27 (
    .O(x15_y27),
    .I0(x13_y25),
    .I1(x12_y28),
    .I2(1'b0),
    .I3(x12_y29)
);

(* keep, dont_touch *)
(* LOC = "X16/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001100001111)
) lut_16_27 (
    .O(x16_y27),
    .I0(x13_y22),
    .I1(x13_y25),
    .I2(x13_y24),
    .I3(x14_y32)
);

(* keep, dont_touch *)
(* LOC = "X17/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100010001011)
) lut_17_27 (
    .O(x17_y27),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x15_y25),
    .I3(x15_y32)
);

(* keep, dont_touch *)
(* LOC = "X18/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010010000101)
) lut_18_27 (
    .O(x18_y27),
    .I0(1'b0),
    .I1(x16_y30),
    .I2(x15_y22),
    .I3(x16_y29)
);

(* keep, dont_touch *)
(* LOC = "X19/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111000100111)
) lut_19_27 (
    .O(x19_y27),
    .I0(1'b0),
    .I1(x16_y22),
    .I2(x16_y27),
    .I3(x17_y27)
);

(* keep, dont_touch *)
(* LOC = "X20/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011000010101)
) lut_20_27 (
    .O(x20_y27),
    .I0(x17_y23),
    .I1(1'b0),
    .I2(x17_y32),
    .I3(x18_y24)
);

(* keep, dont_touch *)
(* LOC = "X21/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100010110011)
) lut_21_27 (
    .O(x21_y27),
    .I0(x18_y22),
    .I1(x19_y23),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X22/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111010100001)
) lut_22_27 (
    .O(x22_y27),
    .I0(1'b0),
    .I1(x19_y29),
    .I2(x20_y25),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X23/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111001111101)
) lut_23_27 (
    .O(x23_y27),
    .I0(x20_y22),
    .I1(x21_y31),
    .I2(x20_y26),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X24/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001000101101)
) lut_24_27 (
    .O(x24_y27),
    .I0(x21_y24),
    .I1(x22_y30),
    .I2(x21_y32),
    .I3(x22_y28)
);

(* keep, dont_touch *)
(* LOC = "X25/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011110110101)
) lut_25_27 (
    .O(x25_y27),
    .I0(x22_y24),
    .I1(x23_y31),
    .I2(x22_y32),
    .I3(x23_y30)
);

(* keep, dont_touch *)
(* LOC = "X26/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111011111101)
) lut_26_27 (
    .O(x26_y27),
    .I0(x23_y25),
    .I1(x24_y28),
    .I2(1'b0),
    .I3(x24_y30)
);

(* keep, dont_touch *)
(* LOC = "X27/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001101000001)
) lut_27_27 (
    .O(x27_y27),
    .I0(x24_y24),
    .I1(x25_y31),
    .I2(x25_y25),
    .I3(x25_y24)
);

(* keep, dont_touch *)
(* LOC = "X28/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000101100011)
) lut_28_27 (
    .O(x28_y27),
    .I0(1'b0),
    .I1(x26_y22),
    .I2(1'b0),
    .I3(x26_y30)
);

(* keep, dont_touch *)
(* LOC = "X29/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110101110100)
) lut_29_27 (
    .O(x29_y27),
    .I0(x27_y23),
    .I1(x26_y30),
    .I2(x27_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X30/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011110111111)
) lut_30_27 (
    .O(x30_y27),
    .I0(1'b0),
    .I1(x28_y30),
    .I2(x27_y32),
    .I3(x27_y28)
);

(* keep, dont_touch *)
(* LOC = "X31/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100111001111)
) lut_31_27 (
    .O(x31_y27),
    .I0(x28_y24),
    .I1(x29_y22),
    .I2(1'b0),
    .I3(x28_y25)
);

(* keep, dont_touch *)
(* LOC = "X32/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110011000011)
) lut_32_27 (
    .O(x32_y27),
    .I0(x30_y26),
    .I1(x30_y22),
    .I2(1'b0),
    .I3(x30_y22)
);

(* keep, dont_touch *)
(* LOC = "X33/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000001000000)
) lut_33_27 (
    .O(x33_y27),
    .I0(1'b0),
    .I1(x30_y23),
    .I2(x31_y28),
    .I3(x31_y28)
);

(* keep, dont_touch *)
(* LOC = "X34/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001111000101)
) lut_34_27 (
    .O(x34_y27),
    .I0(x32_y26),
    .I1(x31_y32),
    .I2(1'b0),
    .I3(x32_y27)
);

(* keep, dont_touch *)
(* LOC = "X35/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101001000000)
) lut_35_27 (
    .O(x35_y27),
    .I0(x33_y26),
    .I1(x33_y25),
    .I2(x32_y24),
    .I3(x33_y24)
);

(* keep, dont_touch *)
(* LOC = "X36/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011101101000)
) lut_36_27 (
    .O(x36_y27),
    .I0(1'b0),
    .I1(x33_y31),
    .I2(1'b0),
    .I3(x33_y25)
);

(* keep, dont_touch *)
(* LOC = "X37/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001010111111)
) lut_37_27 (
    .O(x37_y27),
    .I0(x34_y23),
    .I1(x35_y30),
    .I2(x35_y22),
    .I3(x35_y28)
);

(* keep, dont_touch *)
(* LOC = "X38/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100000100010)
) lut_38_27 (
    .O(x38_y27),
    .I0(x36_y23),
    .I1(x35_y28),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X39/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011101101001)
) lut_39_27 (
    .O(x39_y27),
    .I0(1'b0),
    .I1(x36_y28),
    .I2(x37_y28),
    .I3(x37_y22)
);

(* keep, dont_touch *)
(* LOC = "X40/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110110101110)
) lut_40_27 (
    .O(x40_y27),
    .I0(1'b0),
    .I1(x37_y30),
    .I2(x38_y23),
    .I3(x38_y28)
);

(* keep, dont_touch *)
(* LOC = "X41/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100000111100)
) lut_41_27 (
    .O(x41_y27),
    .I0(x39_y25),
    .I1(1'b0),
    .I2(x38_y27),
    .I3(x39_y27)
);

(* keep, dont_touch *)
(* LOC = "X42/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010100101011)
) lut_42_27 (
    .O(x42_y27),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x40_y25),
    .I3(x40_y27)
);

(* keep, dont_touch *)
(* LOC = "X43/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111101110100)
) lut_43_27 (
    .O(x43_y27),
    .I0(x41_y23),
    .I1(x41_y25),
    .I2(x41_y23),
    .I3(x41_y32)
);

(* keep, dont_touch *)
(* LOC = "X44/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010010100110)
) lut_44_27 (
    .O(x44_y27),
    .I0(1'b0),
    .I1(x41_y29),
    .I2(x42_y24),
    .I3(x42_y24)
);

(* keep, dont_touch *)
(* LOC = "X45/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110110001111)
) lut_45_27 (
    .O(x45_y27),
    .I0(x42_y27),
    .I1(x42_y24),
    .I2(x43_y32),
    .I3(x43_y29)
);

(* keep, dont_touch *)
(* LOC = "X46/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011010101100)
) lut_46_27 (
    .O(x46_y27),
    .I0(x44_y22),
    .I1(1'b0),
    .I2(x44_y24),
    .I3(x43_y27)
);

(* keep, dont_touch *)
(* LOC = "X47/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101110000000)
) lut_47_27 (
    .O(x47_y27),
    .I0(x45_y31),
    .I1(1'b0),
    .I2(x44_y23),
    .I3(x44_y30)
);

(* keep, dont_touch *)
(* LOC = "X48/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010100110100)
) lut_48_27 (
    .O(x48_y27),
    .I0(x46_y24),
    .I1(x45_y26),
    .I2(x45_y30),
    .I3(x46_y22)
);

(* keep, dont_touch *)
(* LOC = "X49/Y27" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110111101010)
) lut_49_27 (
    .O(x49_y27),
    .I0(x46_y31),
    .I1(x47_y27),
    .I2(1'b0),
    .I3(x46_y23)
);

(* keep, dont_touch *)
(* LOC = "X0/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111101000000)
) lut_0_28 (
    .O(x0_y28),
    .I0(in7),
    .I1(1'b0),
    .I2(in4),
    .I3(in5)
);

(* keep, dont_touch *)
(* LOC = "X1/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010111100111)
) lut_1_28 (
    .O(x1_y28),
    .I0(1'b0),
    .I1(in3),
    .I2(in9),
    .I3(in6)
);

(* keep, dont_touch *)
(* LOC = "X2/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101101011010)
) lut_2_28 (
    .O(x2_y28),
    .I0(in8),
    .I1(in3),
    .I2(1'b0),
    .I3(in9)
);

(* keep, dont_touch *)
(* LOC = "X3/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010010001011)
) lut_3_28 (
    .O(x3_y28),
    .I0(x1_y33),
    .I1(in9),
    .I2(x1_y33),
    .I3(in2)
);

(* keep, dont_touch *)
(* LOC = "X4/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100000000010)
) lut_4_28 (
    .O(x4_y28),
    .I0(x2_y24),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x2_y26)
);

(* keep, dont_touch *)
(* LOC = "X5/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111101010010)
) lut_5_28 (
    .O(x5_y28),
    .I0(x2_y26),
    .I1(1'b0),
    .I2(x3_y23),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X6/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011010000001)
) lut_6_28 (
    .O(x6_y28),
    .I0(x3_y30),
    .I1(x4_y25),
    .I2(1'b0),
    .I3(x3_y32)
);

(* keep, dont_touch *)
(* LOC = "X7/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100000100000)
) lut_7_28 (
    .O(x7_y28),
    .I0(x5_y27),
    .I1(x5_y32),
    .I2(x5_y24),
    .I3(x4_y25)
);

(* keep, dont_touch *)
(* LOC = "X8/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001010101001)
) lut_8_28 (
    .O(x8_y28),
    .I0(x5_y28),
    .I1(x6_y29),
    .I2(x5_y25),
    .I3(x5_y25)
);

(* keep, dont_touch *)
(* LOC = "X9/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111101111010)
) lut_9_28 (
    .O(x9_y28),
    .I0(1'b0),
    .I1(x6_y27),
    .I2(x5_y25),
    .I3(x5_y25)
);

(* keep, dont_touch *)
(* LOC = "X10/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110110001111)
) lut_10_28 (
    .O(x10_y28),
    .I0(x8_y26),
    .I1(x7_y24),
    .I2(x7_y27),
    .I3(x7_y27)
);

(* keep, dont_touch *)
(* LOC = "X11/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001010001111)
) lut_11_28 (
    .O(x11_y28),
    .I0(x9_y26),
    .I1(x8_y23),
    .I2(1'b0),
    .I3(x9_y27)
);

(* keep, dont_touch *)
(* LOC = "X12/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110011010100)
) lut_12_28 (
    .O(x12_y28),
    .I0(x9_y29),
    .I1(x10_y32),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X13/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100001110000)
) lut_13_28 (
    .O(x13_y28),
    .I0(x10_y30),
    .I1(1'b0),
    .I2(x10_y25),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X14/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110000001101)
) lut_14_28 (
    .O(x14_y28),
    .I0(1'b0),
    .I1(x12_y24),
    .I2(x11_y24),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X15/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110100101010)
) lut_15_28 (
    .O(x15_y28),
    .I0(x13_y32),
    .I1(x13_y32),
    .I2(1'b0),
    .I3(x13_y26)
);

(* keep, dont_touch *)
(* LOC = "X16/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010111101011)
) lut_16_28 (
    .O(x16_y28),
    .I0(x13_y28),
    .I1(1'b0),
    .I2(x13_y30),
    .I3(x14_y28)
);

(* keep, dont_touch *)
(* LOC = "X17/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110110000101)
) lut_17_28 (
    .O(x17_y28),
    .I0(x14_y26),
    .I1(x15_y33),
    .I2(x14_y23),
    .I3(x15_y27)
);

(* keep, dont_touch *)
(* LOC = "X18/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101111000010)
) lut_18_28 (
    .O(x18_y28),
    .I0(x15_y25),
    .I1(x15_y26),
    .I2(x16_y27),
    .I3(x16_y29)
);

(* keep, dont_touch *)
(* LOC = "X19/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001101101011)
) lut_19_28 (
    .O(x19_y28),
    .I0(1'b0),
    .I1(x16_y25),
    .I2(1'b0),
    .I3(x17_y33)
);

(* keep, dont_touch *)
(* LOC = "X20/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011110010111)
) lut_20_28 (
    .O(x20_y28),
    .I0(x17_y25),
    .I1(x17_y24),
    .I2(x18_y31),
    .I3(x18_y27)
);

(* keep, dont_touch *)
(* LOC = "X21/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111010101111)
) lut_21_28 (
    .O(x21_y28),
    .I0(x18_y28),
    .I1(x18_y26),
    .I2(x19_y33),
    .I3(x18_y32)
);

(* keep, dont_touch *)
(* LOC = "X22/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001111110010)
) lut_22_28 (
    .O(x22_y28),
    .I0(x20_y32),
    .I1(1'b0),
    .I2(x19_y27),
    .I3(x20_y24)
);

(* keep, dont_touch *)
(* LOC = "X23/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000100000111)
) lut_23_28 (
    .O(x23_y28),
    .I0(x21_y30),
    .I1(1'b0),
    .I2(x21_y31),
    .I3(x21_y23)
);

(* keep, dont_touch *)
(* LOC = "X24/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000001110110)
) lut_24_28 (
    .O(x24_y28),
    .I0(1'b0),
    .I1(x22_y26),
    .I2(1'b0),
    .I3(x22_y23)
);

(* keep, dont_touch *)
(* LOC = "X25/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101001010110)
) lut_25_28 (
    .O(x25_y28),
    .I0(x23_y28),
    .I1(1'b0),
    .I2(x23_y28),
    .I3(x23_y23)
);

(* keep, dont_touch *)
(* LOC = "X26/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110000011011)
) lut_26_28 (
    .O(x26_y28),
    .I0(1'b0),
    .I1(x23_y32),
    .I2(x23_y26),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X27/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111011011110)
) lut_27_28 (
    .O(x27_y28),
    .I0(x24_y27),
    .I1(x24_y31),
    .I2(1'b0),
    .I3(x25_y24)
);

(* keep, dont_touch *)
(* LOC = "X28/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001001000001)
) lut_28_28 (
    .O(x28_y28),
    .I0(x26_y31),
    .I1(1'b0),
    .I2(x25_y23),
    .I3(x25_y27)
);

(* keep, dont_touch *)
(* LOC = "X29/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111101010110)
) lut_29_28 (
    .O(x29_y28),
    .I0(1'b0),
    .I1(x27_y33),
    .I2(x27_y30),
    .I3(x26_y26)
);

(* keep, dont_touch *)
(* LOC = "X30/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100111010111)
) lut_30_28 (
    .O(x30_y28),
    .I0(x27_y24),
    .I1(x28_y26),
    .I2(x27_y31),
    .I3(x27_y23)
);

(* keep, dont_touch *)
(* LOC = "X31/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111011110110)
) lut_31_28 (
    .O(x31_y28),
    .I0(x28_y33),
    .I1(x28_y25),
    .I2(x29_y31),
    .I3(x29_y31)
);

(* keep, dont_touch *)
(* LOC = "X32/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100101010111)
) lut_32_28 (
    .O(x32_y28),
    .I0(1'b0),
    .I1(x29_y31),
    .I2(x29_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X33/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100010101111)
) lut_33_28 (
    .O(x33_y28),
    .I0(x31_y26),
    .I1(x31_y29),
    .I2(x31_y31),
    .I3(x31_y28)
);

(* keep, dont_touch *)
(* LOC = "X34/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011000011010)
) lut_34_28 (
    .O(x34_y28),
    .I0(x31_y23),
    .I1(x31_y24),
    .I2(x31_y31),
    .I3(x32_y24)
);

(* keep, dont_touch *)
(* LOC = "X35/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000110001111)
) lut_35_28 (
    .O(x35_y28),
    .I0(x33_y25),
    .I1(1'b0),
    .I2(x33_y31),
    .I3(x32_y33)
);

(* keep, dont_touch *)
(* LOC = "X36/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000101000100)
) lut_36_28 (
    .O(x36_y28),
    .I0(x34_y33),
    .I1(x33_y29),
    .I2(1'b0),
    .I3(x33_y29)
);

(* keep, dont_touch *)
(* LOC = "X37/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111111001101)
) lut_37_28 (
    .O(x37_y28),
    .I0(x34_y28),
    .I1(x34_y33),
    .I2(1'b0),
    .I3(x35_y31)
);

(* keep, dont_touch *)
(* LOC = "X38/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011100100011)
) lut_38_28 (
    .O(x38_y28),
    .I0(x35_y31),
    .I1(x35_y27),
    .I2(x36_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X39/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010101100100)
) lut_39_28 (
    .O(x39_y28),
    .I0(x36_y25),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x36_y23)
);

(* keep, dont_touch *)
(* LOC = "X40/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111110000001)
) lut_40_28 (
    .O(x40_y28),
    .I0(x37_y28),
    .I1(x38_y25),
    .I2(x38_y24),
    .I3(x37_y23)
);

(* keep, dont_touch *)
(* LOC = "X41/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011010111100)
) lut_41_28 (
    .O(x41_y28),
    .I0(x38_y27),
    .I1(x38_y27),
    .I2(x38_y25),
    .I3(x39_y25)
);

(* keep, dont_touch *)
(* LOC = "X42/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011110011011)
) lut_42_28 (
    .O(x42_y28),
    .I0(x39_y32),
    .I1(x40_y23),
    .I2(1'b0),
    .I3(x39_y25)
);

(* keep, dont_touch *)
(* LOC = "X43/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011100010010)
) lut_43_28 (
    .O(x43_y28),
    .I0(x41_y31),
    .I1(x40_y24),
    .I2(1'b0),
    .I3(x41_y29)
);

(* keep, dont_touch *)
(* LOC = "X44/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111100101110)
) lut_44_28 (
    .O(x44_y28),
    .I0(x41_y31),
    .I1(x42_y27),
    .I2(x41_y33),
    .I3(x41_y23)
);

(* keep, dont_touch *)
(* LOC = "X45/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011100000000)
) lut_45_28 (
    .O(x45_y28),
    .I0(x43_y33),
    .I1(x42_y29),
    .I2(x42_y24),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X46/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010101010000)
) lut_46_28 (
    .O(x46_y28),
    .I0(x43_y27),
    .I1(x43_y27),
    .I2(x44_y26),
    .I3(x43_y31)
);

(* keep, dont_touch *)
(* LOC = "X47/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110101110100)
) lut_47_28 (
    .O(x47_y28),
    .I0(x45_y29),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x44_y28)
);

(* keep, dont_touch *)
(* LOC = "X48/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110010110010)
) lut_48_28 (
    .O(x48_y28),
    .I0(1'b0),
    .I1(x46_y32),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X49/Y28" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110000100111)
) lut_49_28 (
    .O(x49_y28),
    .I0(x46_y24),
    .I1(x46_y28),
    .I2(x47_y24),
    .I3(x46_y31)
);

(* keep, dont_touch *)
(* LOC = "X0/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111010111001)
) lut_0_29 (
    .O(x0_y29),
    .I0(1'b0),
    .I1(in9),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X1/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000001000000)
) lut_1_29 (
    .O(x1_y29),
    .I0(1'b0),
    .I1(in7),
    .I2(in1),
    .I3(in1)
);

(* keep, dont_touch *)
(* LOC = "X2/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111111000101)
) lut_2_29 (
    .O(x2_y29),
    .I0(1'b0),
    .I1(in2),
    .I2(1'b0),
    .I3(in4)
);

(* keep, dont_touch *)
(* LOC = "X3/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011111001000)
) lut_3_29 (
    .O(x3_y29),
    .I0(1'b0),
    .I1(x1_y30),
    .I2(in4),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X4/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011001100000)
) lut_4_29 (
    .O(x4_y29),
    .I0(1'b0),
    .I1(x2_y34),
    .I2(1'b0),
    .I3(x1_y33)
);

(* keep, dont_touch *)
(* LOC = "X5/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011001000010)
) lut_5_29 (
    .O(x5_y29),
    .I0(1'b0),
    .I1(x2_y30),
    .I2(x2_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X6/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011110110001)
) lut_6_29 (
    .O(x6_y29),
    .I0(1'b0),
    .I1(x4_y31),
    .I2(x3_y29),
    .I3(x4_y24)
);

(* keep, dont_touch *)
(* LOC = "X7/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011101101011)
) lut_7_29 (
    .O(x7_y29),
    .I0(x5_y28),
    .I1(x5_y27),
    .I2(1'b0),
    .I3(x5_y34)
);

(* keep, dont_touch *)
(* LOC = "X8/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100000110011)
) lut_8_29 (
    .O(x8_y29),
    .I0(x5_y28),
    .I1(x5_y29),
    .I2(x6_y27),
    .I3(x6_y32)
);

(* keep, dont_touch *)
(* LOC = "X9/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111111001000)
) lut_9_29 (
    .O(x9_y29),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x6_y27),
    .I3(x6_y32)
);

(* keep, dont_touch *)
(* LOC = "X10/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011000011100)
) lut_10_29 (
    .O(x10_y29),
    .I0(x8_y31),
    .I1(1'b0),
    .I2(x7_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X11/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111110010011)
) lut_11_29 (
    .O(x11_y29),
    .I0(x8_y34),
    .I1(x8_y25),
    .I2(x9_y30),
    .I3(x9_y27)
);

(* keep, dont_touch *)
(* LOC = "X12/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001010101000)
) lut_12_29 (
    .O(x12_y29),
    .I0(1'b0),
    .I1(x9_y25),
    .I2(x10_y25),
    .I3(x9_y28)
);

(* keep, dont_touch *)
(* LOC = "X13/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101110001001)
) lut_13_29 (
    .O(x13_y29),
    .I0(x10_y31),
    .I1(x11_y33),
    .I2(x11_y26),
    .I3(x11_y25)
);

(* keep, dont_touch *)
(* LOC = "X14/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001100101110)
) lut_14_29 (
    .O(x14_y29),
    .I0(x12_y25),
    .I1(1'b0),
    .I2(x12_y25),
    .I3(x12_y33)
);

(* keep, dont_touch *)
(* LOC = "X15/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001011101000)
) lut_15_29 (
    .O(x15_y29),
    .I0(x12_y27),
    .I1(x12_y30),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X16/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001010011111)
) lut_16_29 (
    .O(x16_y29),
    .I0(x14_y29),
    .I1(x14_y24),
    .I2(x13_y24),
    .I3(x13_y31)
);

(* keep, dont_touch *)
(* LOC = "X17/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001111011001)
) lut_17_29 (
    .O(x17_y29),
    .I0(x15_y31),
    .I1(x15_y33),
    .I2(x14_y30),
    .I3(x14_y28)
);

(* keep, dont_touch *)
(* LOC = "X18/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011001010000)
) lut_18_29 (
    .O(x18_y29),
    .I0(x16_y26),
    .I1(x16_y30),
    .I2(x15_y25),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X19/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110000101100)
) lut_19_29 (
    .O(x19_y29),
    .I0(x17_y33),
    .I1(x17_y24),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X20/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100010001010)
) lut_20_29 (
    .O(x20_y29),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x18_y29)
);

(* keep, dont_touch *)
(* LOC = "X21/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010100110100)
) lut_21_29 (
    .O(x21_y29),
    .I0(x18_y34),
    .I1(x19_y30),
    .I2(x19_y24),
    .I3(x18_y32)
);

(* keep, dont_touch *)
(* LOC = "X22/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100100111000)
) lut_22_29 (
    .O(x22_y29),
    .I0(x20_y27),
    .I1(x20_y28),
    .I2(x19_y24),
    .I3(x19_y24)
);

(* keep, dont_touch *)
(* LOC = "X23/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001001111001)
) lut_23_29 (
    .O(x23_y29),
    .I0(x21_y28),
    .I1(x20_y24),
    .I2(1'b0),
    .I3(x20_y33)
);

(* keep, dont_touch *)
(* LOC = "X24/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111111001011)
) lut_24_29 (
    .O(x24_y29),
    .I0(x21_y28),
    .I1(x22_y26),
    .I2(x22_y29),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X25/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011001110111)
) lut_25_29 (
    .O(x25_y29),
    .I0(1'b0),
    .I1(x23_y27),
    .I2(x22_y34),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X26/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111000000101)
) lut_26_29 (
    .O(x26_y29),
    .I0(x23_y33),
    .I1(1'b0),
    .I2(x23_y29),
    .I3(x24_y27)
);

(* keep, dont_touch *)
(* LOC = "X27/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110000011110)
) lut_27_29 (
    .O(x27_y29),
    .I0(x24_y32),
    .I1(x24_y25),
    .I2(x24_y31),
    .I3(x25_y34)
);

(* keep, dont_touch *)
(* LOC = "X28/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010011111011)
) lut_28_29 (
    .O(x28_y29),
    .I0(x25_y32),
    .I1(1'b0),
    .I2(x25_y30),
    .I3(x25_y25)
);

(* keep, dont_touch *)
(* LOC = "X29/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010111001000)
) lut_29_29 (
    .O(x29_y29),
    .I0(1'b0),
    .I1(x27_y27),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X30/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101001101110)
) lut_30_29 (
    .O(x30_y29),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x27_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X31/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101011100001)
) lut_31_29 (
    .O(x31_y29),
    .I0(1'b0),
    .I1(x29_y27),
    .I2(x28_y31),
    .I3(x29_y25)
);

(* keep, dont_touch *)
(* LOC = "X32/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000100010011)
) lut_32_29 (
    .O(x32_y29),
    .I0(x30_y31),
    .I1(1'b0),
    .I2(x29_y33),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X33/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000011010110)
) lut_33_29 (
    .O(x33_y29),
    .I0(x31_y34),
    .I1(x30_y33),
    .I2(x30_y31),
    .I3(x31_y27)
);

(* keep, dont_touch *)
(* LOC = "X34/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000001000001)
) lut_34_29 (
    .O(x34_y29),
    .I0(x32_y27),
    .I1(x32_y28),
    .I2(x31_y27),
    .I3(x31_y29)
);

(* keep, dont_touch *)
(* LOC = "X35/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000011001010)
) lut_35_29 (
    .O(x35_y29),
    .I0(x32_y28),
    .I1(x33_y31),
    .I2(1'b0),
    .I3(x32_y25)
);

(* keep, dont_touch *)
(* LOC = "X36/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010000100000)
) lut_36_29 (
    .O(x36_y29),
    .I0(x33_y26),
    .I1(x34_y32),
    .I2(x34_y24),
    .I3(x33_y34)
);

(* keep, dont_touch *)
(* LOC = "X37/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111100011110)
) lut_37_29 (
    .O(x37_y29),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x34_y29),
    .I3(x34_y29)
);

(* keep, dont_touch *)
(* LOC = "X38/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110111000011)
) lut_38_29 (
    .O(x38_y29),
    .I0(x36_y25),
    .I1(1'b0),
    .I2(x36_y26),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X39/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010101001110)
) lut_39_29 (
    .O(x39_y29),
    .I0(x37_y34),
    .I1(x37_y24),
    .I2(x36_y24),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X40/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100000100101)
) lut_40_29 (
    .O(x40_y29),
    .I0(1'b0),
    .I1(x38_y29),
    .I2(1'b0),
    .I3(x38_y27)
);

(* keep, dont_touch *)
(* LOC = "X41/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100001010100)
) lut_41_29 (
    .O(x41_y29),
    .I0(x39_y30),
    .I1(x39_y27),
    .I2(x39_y25),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X42/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001001111001)
) lut_42_29 (
    .O(x42_y29),
    .I0(x40_y30),
    .I1(x40_y30),
    .I2(1'b0),
    .I3(x39_y26)
);

(* keep, dont_touch *)
(* LOC = "X43/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011111101110)
) lut_43_29 (
    .O(x43_y29),
    .I0(x40_y26),
    .I1(1'b0),
    .I2(x41_y33),
    .I3(x41_y27)
);

(* keep, dont_touch *)
(* LOC = "X44/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110111010000)
) lut_44_29 (
    .O(x44_y29),
    .I0(x41_y28),
    .I1(x41_y31),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X45/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000010101110)
) lut_45_29 (
    .O(x45_y29),
    .I0(x43_y31),
    .I1(x43_y27),
    .I2(1'b0),
    .I3(x42_y31)
);

(* keep, dont_touch *)
(* LOC = "X46/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000100100110)
) lut_46_29 (
    .O(x46_y29),
    .I0(x44_y33),
    .I1(x44_y27),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X47/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010011010111)
) lut_47_29 (
    .O(x47_y29),
    .I0(x45_y32),
    .I1(1'b0),
    .I2(x44_y30),
    .I3(x45_y28)
);

(* keep, dont_touch *)
(* LOC = "X48/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110100000100)
) lut_48_29 (
    .O(x48_y29),
    .I0(x46_y24),
    .I1(x46_y27),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X49/Y29" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100001000100)
) lut_49_29 (
    .O(x49_y29),
    .I0(x47_y34),
    .I1(x47_y34),
    .I2(x46_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X0/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000111111101)
) lut_0_30 (
    .O(x0_y30),
    .I0(in3),
    .I1(in0),
    .I2(in9),
    .I3(in9)
);

(* keep, dont_touch *)
(* LOC = "X1/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001111000001)
) lut_1_30 (
    .O(x1_y30),
    .I0(in2),
    .I1(in5),
    .I2(1'b0),
    .I3(in1)
);

(* keep, dont_touch *)
(* LOC = "X2/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110110110101)
) lut_2_30 (
    .O(x2_y30),
    .I0(in9),
    .I1(1'b0),
    .I2(in9),
    .I3(in8)
);

(* keep, dont_touch *)
(* LOC = "X3/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011111100101)
) lut_3_30 (
    .O(x3_y30),
    .I0(in9),
    .I1(x1_y28),
    .I2(in4),
    .I3(x1_y32)
);

(* keep, dont_touch *)
(* LOC = "X4/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111010110101)
) lut_4_30 (
    .O(x4_y30),
    .I0(x2_y32),
    .I1(x1_y32),
    .I2(x2_y33),
    .I3(x1_y33)
);

(* keep, dont_touch *)
(* LOC = "X5/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100010000001)
) lut_5_30 (
    .O(x5_y30),
    .I0(x2_y31),
    .I1(x3_y31),
    .I2(x2_y35),
    .I3(x3_y26)
);

(* keep, dont_touch *)
(* LOC = "X6/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100010011100)
) lut_6_30 (
    .O(x6_y30),
    .I0(x3_y25),
    .I1(1'b0),
    .I2(x4_y27),
    .I3(x4_y27)
);

(* keep, dont_touch *)
(* LOC = "X7/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101100011011)
) lut_7_30 (
    .O(x7_y30),
    .I0(1'b0),
    .I1(x5_y33),
    .I2(x4_y27),
    .I3(x5_y26)
);

(* keep, dont_touch *)
(* LOC = "X8/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111111011000)
) lut_8_30 (
    .O(x8_y30),
    .I0(x6_y33),
    .I1(x6_y25),
    .I2(1'b0),
    .I3(x5_y30)
);

(* keep, dont_touch *)
(* LOC = "X9/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101110110001)
) lut_9_30 (
    .O(x9_y30),
    .I0(x6_y29),
    .I1(x6_y30),
    .I2(1'b0),
    .I3(x5_y30)
);

(* keep, dont_touch *)
(* LOC = "X10/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110110101001)
) lut_10_30 (
    .O(x10_y30),
    .I0(1'b0),
    .I1(x8_y27),
    .I2(x8_y32),
    .I3(x8_y32)
);

(* keep, dont_touch *)
(* LOC = "X11/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101111101100)
) lut_11_30 (
    .O(x11_y30),
    .I0(1'b0),
    .I1(x8_y31),
    .I2(x8_y29),
    .I3(x8_y29)
);

(* keep, dont_touch *)
(* LOC = "X12/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001101001101)
) lut_12_30 (
    .O(x12_y30),
    .I0(1'b0),
    .I1(x9_y26),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X13/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011010011100)
) lut_13_30 (
    .O(x13_y30),
    .I0(x11_y29),
    .I1(x11_y34),
    .I2(x11_y31),
    .I3(x10_y31)
);

(* keep, dont_touch *)
(* LOC = "X14/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100110000010)
) lut_14_30 (
    .O(x14_y30),
    .I0(x12_y34),
    .I1(x11_y30),
    .I2(x12_y29),
    .I3(x12_y33)
);

(* keep, dont_touch *)
(* LOC = "X15/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100110111110)
) lut_15_30 (
    .O(x15_y30),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x12_y25)
);

(* keep, dont_touch *)
(* LOC = "X16/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100011101111)
) lut_16_30 (
    .O(x16_y30),
    .I0(x13_y34),
    .I1(1'b0),
    .I2(x13_y31),
    .I3(x13_y26)
);

(* keep, dont_touch *)
(* LOC = "X17/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001110010011)
) lut_17_30 (
    .O(x17_y30),
    .I0(x15_y26),
    .I1(x14_y25),
    .I2(x15_y26),
    .I3(x15_y30)
);

(* keep, dont_touch *)
(* LOC = "X18/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101101010111)
) lut_18_30 (
    .O(x18_y30),
    .I0(x16_y28),
    .I1(x15_y34),
    .I2(x16_y25),
    .I3(x15_y30)
);

(* keep, dont_touch *)
(* LOC = "X19/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011011101001)
) lut_19_30 (
    .O(x19_y30),
    .I0(1'b0),
    .I1(x17_y28),
    .I2(x16_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X20/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110101010010)
) lut_20_30 (
    .O(x20_y30),
    .I0(x17_y33),
    .I1(x17_y29),
    .I2(x18_y29),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X21/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101001111010)
) lut_21_30 (
    .O(x21_y30),
    .I0(x18_y26),
    .I1(x19_y25),
    .I2(x18_y27),
    .I3(x18_y35)
);

(* keep, dont_touch *)
(* LOC = "X22/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101101010001)
) lut_22_30 (
    .O(x22_y30),
    .I0(x19_y30),
    .I1(x19_y30),
    .I2(1'b0),
    .I3(x20_y34)
);

(* keep, dont_touch *)
(* LOC = "X23/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001111000100)
) lut_23_30 (
    .O(x23_y30),
    .I0(x20_y25),
    .I1(x20_y35),
    .I2(x20_y29),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X24/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001110010010)
) lut_24_30 (
    .O(x24_y30),
    .I0(x21_y30),
    .I1(x21_y35),
    .I2(x22_y35),
    .I3(x22_y25)
);

(* keep, dont_touch *)
(* LOC = "X25/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010001000000)
) lut_25_30 (
    .O(x25_y30),
    .I0(x23_y30),
    .I1(x23_y32),
    .I2(1'b0),
    .I3(x22_y27)
);

(* keep, dont_touch *)
(* LOC = "X26/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001000101001)
) lut_26_30 (
    .O(x26_y30),
    .I0(1'b0),
    .I1(x24_y30),
    .I2(x23_y34),
    .I3(x24_y27)
);

(* keep, dont_touch *)
(* LOC = "X27/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111111101010)
) lut_27_30 (
    .O(x27_y30),
    .I0(x24_y34),
    .I1(x25_y25),
    .I2(x25_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X28/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001010010010)
) lut_28_30 (
    .O(x28_y30),
    .I0(x25_y27),
    .I1(x26_y26),
    .I2(x25_y30),
    .I3(x25_y29)
);

(* keep, dont_touch *)
(* LOC = "X29/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110111100011)
) lut_29_30 (
    .O(x29_y30),
    .I0(x27_y27),
    .I1(x26_y35),
    .I2(x27_y35),
    .I3(x26_y33)
);

(* keep, dont_touch *)
(* LOC = "X30/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101011100101)
) lut_30_30 (
    .O(x30_y30),
    .I0(x27_y25),
    .I1(x27_y25),
    .I2(x27_y25),
    .I3(x28_y26)
);

(* keep, dont_touch *)
(* LOC = "X31/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010000110100)
) lut_31_30 (
    .O(x31_y30),
    .I0(x28_y33),
    .I1(x28_y28),
    .I2(x29_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X32/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100001000010)
) lut_32_30 (
    .O(x32_y30),
    .I0(1'b0),
    .I1(x30_y35),
    .I2(x29_y33),
    .I3(x29_y35)
);

(* keep, dont_touch *)
(* LOC = "X33/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011000011100)
) lut_33_30 (
    .O(x33_y30),
    .I0(x31_y34),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X34/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100010000000)
) lut_34_30 (
    .O(x34_y30),
    .I0(x32_y26),
    .I1(x32_y32),
    .I2(1'b0),
    .I3(x32_y30)
);

(* keep, dont_touch *)
(* LOC = "X35/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111111011110)
) lut_35_30 (
    .O(x35_y30),
    .I0(x33_y31),
    .I1(1'b0),
    .I2(x32_y35),
    .I3(x33_y27)
);

(* keep, dont_touch *)
(* LOC = "X36/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000110001000)
) lut_36_30 (
    .O(x36_y30),
    .I0(x33_y35),
    .I1(x34_y28),
    .I2(x34_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X37/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001100100101)
) lut_37_30 (
    .O(x37_y30),
    .I0(x34_y27),
    .I1(x35_y29),
    .I2(x35_y34),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X38/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000101001100)
) lut_38_30 (
    .O(x38_y30),
    .I0(x35_y31),
    .I1(x35_y28),
    .I2(x35_y33),
    .I3(x35_y26)
);

(* keep, dont_touch *)
(* LOC = "X39/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101011111010)
) lut_39_30 (
    .O(x39_y30),
    .I0(1'b0),
    .I1(x37_y33),
    .I2(1'b0),
    .I3(x37_y25)
);

(* keep, dont_touch *)
(* LOC = "X40/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000100101101)
) lut_40_30 (
    .O(x40_y30),
    .I0(x37_y33),
    .I1(x38_y27),
    .I2(x38_y29),
    .I3(x37_y27)
);

(* keep, dont_touch *)
(* LOC = "X41/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001001100111)
) lut_41_30 (
    .O(x41_y30),
    .I0(x38_y31),
    .I1(1'b0),
    .I2(x39_y32),
    .I3(x39_y34)
);

(* keep, dont_touch *)
(* LOC = "X42/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101011111001)
) lut_42_30 (
    .O(x42_y30),
    .I0(x40_y28),
    .I1(x39_y35),
    .I2(1'b0),
    .I3(x40_y35)
);

(* keep, dont_touch *)
(* LOC = "X43/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000110010111)
) lut_43_30 (
    .O(x43_y30),
    .I0(1'b0),
    .I1(x40_y32),
    .I2(x41_y34),
    .I3(x40_y31)
);

(* keep, dont_touch *)
(* LOC = "X44/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000110110011)
) lut_44_30 (
    .O(x44_y30),
    .I0(x41_y33),
    .I1(x42_y30),
    .I2(1'b0),
    .I3(x42_y29)
);

(* keep, dont_touch *)
(* LOC = "X45/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010110101111)
) lut_45_30 (
    .O(x45_y30),
    .I0(1'b0),
    .I1(x42_y35),
    .I2(x43_y25),
    .I3(x43_y28)
);

(* keep, dont_touch *)
(* LOC = "X46/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010000010000)
) lut_46_30 (
    .O(x46_y30),
    .I0(1'b0),
    .I1(x44_y26),
    .I2(x44_y27),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X47/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001001110000)
) lut_47_30 (
    .O(x47_y30),
    .I0(x44_y29),
    .I1(x44_y28),
    .I2(x44_y26),
    .I3(x45_y34)
);

(* keep, dont_touch *)
(* LOC = "X48/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101111111100)
) lut_48_30 (
    .O(x48_y30),
    .I0(1'b0),
    .I1(x45_y34),
    .I2(x46_y28),
    .I3(x45_y32)
);

(* keep, dont_touch *)
(* LOC = "X49/Y30" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011001111010)
) lut_49_30 (
    .O(x49_y30),
    .I0(x46_y27),
    .I1(x46_y33),
    .I2(1'b0),
    .I3(x47_y31)
);

(* keep, dont_touch *)
(* LOC = "X0/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001111010110)
) lut_0_31 (
    .O(x0_y31),
    .I0(1'b0),
    .I1(in2),
    .I2(in1),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X1/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000001101101)
) lut_1_31 (
    .O(x1_y31),
    .I0(1'b0),
    .I1(1'b0),
    .I2(in8),
    .I3(in6)
);

(* keep, dont_touch *)
(* LOC = "X2/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011100011011)
) lut_2_31 (
    .O(x2_y31),
    .I0(in0),
    .I1(in5),
    .I2(in1),
    .I3(in4)
);

(* keep, dont_touch *)
(* LOC = "X3/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101001000001)
) lut_3_31 (
    .O(x3_y31),
    .I0(in3),
    .I1(in8),
    .I2(x1_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X4/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111000000010)
) lut_4_31 (
    .O(x4_y31),
    .I0(x2_y35),
    .I1(x1_y34),
    .I2(x1_y36),
    .I3(x2_y29)
);

(* keep, dont_touch *)
(* LOC = "X5/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011011111100)
) lut_5_31 (
    .O(x5_y31),
    .I0(1'b0),
    .I1(x2_y33),
    .I2(x2_y36),
    .I3(x3_y36)
);

(* keep, dont_touch *)
(* LOC = "X6/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011111110111)
) lut_6_31 (
    .O(x6_y31),
    .I0(x4_y36),
    .I1(x4_y29),
    .I2(x3_y33),
    .I3(x4_y28)
);

(* keep, dont_touch *)
(* LOC = "X7/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101011000110)
) lut_7_31 (
    .O(x7_y31),
    .I0(x4_y32),
    .I1(x5_y35),
    .I2(x5_y26),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X8/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110000011110)
) lut_8_31 (
    .O(x8_y31),
    .I0(x6_y36),
    .I1(x6_y33),
    .I2(x5_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X9/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001011011100)
) lut_9_31 (
    .O(x9_y31),
    .I0(x7_y27),
    .I1(x6_y35),
    .I2(x5_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X10/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101111110110)
) lut_10_31 (
    .O(x10_y31),
    .I0(x7_y29),
    .I1(1'b0),
    .I2(x8_y30),
    .I3(x7_y29)
);

(* keep, dont_touch *)
(* LOC = "X11/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000111010010)
) lut_11_31 (
    .O(x11_y31),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x9_y31),
    .I3(x9_y29)
);

(* keep, dont_touch *)
(* LOC = "X12/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110010000010)
) lut_12_31 (
    .O(x12_y31),
    .I0(x10_y27),
    .I1(x9_y34),
    .I2(x9_y27),
    .I3(x10_y28)
);

(* keep, dont_touch *)
(* LOC = "X13/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100000011111)
) lut_13_31 (
    .O(x13_y31),
    .I0(x10_y29),
    .I1(x11_y28),
    .I2(x10_y33),
    .I3(x10_y33)
);

(* keep, dont_touch *)
(* LOC = "X14/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000001000101)
) lut_14_31 (
    .O(x14_y31),
    .I0(x12_y32),
    .I1(1'b0),
    .I2(x11_y29),
    .I3(x11_y34)
);

(* keep, dont_touch *)
(* LOC = "X15/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000100010110)
) lut_15_31 (
    .O(x15_y31),
    .I0(x13_y34),
    .I1(1'b0),
    .I2(x12_y31),
    .I3(x12_y33)
);

(* keep, dont_touch *)
(* LOC = "X16/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101010110100)
) lut_16_31 (
    .O(x16_y31),
    .I0(1'b0),
    .I1(x14_y26),
    .I2(x14_y29),
    .I3(x13_y26)
);

(* keep, dont_touch *)
(* LOC = "X17/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000101111101)
) lut_17_31 (
    .O(x17_y31),
    .I0(x14_y36),
    .I1(x15_y31),
    .I2(x15_y31),
    .I3(x15_y28)
);

(* keep, dont_touch *)
(* LOC = "X18/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000110001100)
) lut_18_31 (
    .O(x18_y31),
    .I0(x15_y34),
    .I1(x15_y33),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X19/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001000011000)
) lut_19_31 (
    .O(x19_y31),
    .I0(x17_y28),
    .I1(x17_y27),
    .I2(x16_y28),
    .I3(x17_y26)
);

(* keep, dont_touch *)
(* LOC = "X20/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011000100011)
) lut_20_31 (
    .O(x20_y31),
    .I0(x18_y29),
    .I1(1'b0),
    .I2(x17_y27),
    .I3(x17_y26)
);

(* keep, dont_touch *)
(* LOC = "X21/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011101011010)
) lut_21_31 (
    .O(x21_y31),
    .I0(x19_y28),
    .I1(x19_y33),
    .I2(x19_y31),
    .I3(x19_y34)
);

(* keep, dont_touch *)
(* LOC = "X22/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100010110000)
) lut_22_31 (
    .O(x22_y31),
    .I0(x20_y31),
    .I1(x19_y32),
    .I2(x19_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X23/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000011000110)
) lut_23_31 (
    .O(x23_y31),
    .I0(x20_y30),
    .I1(x21_y32),
    .I2(x20_y33),
    .I3(x21_y32)
);

(* keep, dont_touch *)
(* LOC = "X24/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000100100011)
) lut_24_31 (
    .O(x24_y31),
    .I0(x21_y34),
    .I1(x21_y30),
    .I2(x21_y35),
    .I3(x21_y26)
);

(* keep, dont_touch *)
(* LOC = "X25/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011100010111)
) lut_25_31 (
    .O(x25_y31),
    .I0(x22_y33),
    .I1(x22_y27),
    .I2(x23_y33),
    .I3(x23_y33)
);

(* keep, dont_touch *)
(* LOC = "X26/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011111000111)
) lut_26_31 (
    .O(x26_y31),
    .I0(x23_y35),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X27/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011000000100)
) lut_27_31 (
    .O(x27_y31),
    .I0(x25_y33),
    .I1(x25_y30),
    .I2(x24_y33),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X28/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111001101100)
) lut_28_31 (
    .O(x28_y31),
    .I0(x26_y32),
    .I1(x26_y30),
    .I2(x26_y33),
    .I3(x25_y26)
);

(* keep, dont_touch *)
(* LOC = "X29/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100001110101)
) lut_29_31 (
    .O(x29_y31),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x26_y26),
    .I3(x26_y36)
);

(* keep, dont_touch *)
(* LOC = "X30/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001000100010)
) lut_30_31 (
    .O(x30_y31),
    .I0(x28_y29),
    .I1(1'b0),
    .I2(x28_y36),
    .I3(x28_y27)
);

(* keep, dont_touch *)
(* LOC = "X31/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101010001100)
) lut_31_31 (
    .O(x31_y31),
    .I0(x29_y34),
    .I1(x28_y28),
    .I2(x29_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X32/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111110000010)
) lut_32_31 (
    .O(x32_y31),
    .I0(1'b0),
    .I1(x29_y34),
    .I2(x30_y33),
    .I3(x29_y35)
);

(* keep, dont_touch *)
(* LOC = "X33/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011010010110)
) lut_33_31 (
    .O(x33_y31),
    .I0(x31_y27),
    .I1(1'b0),
    .I2(x30_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X34/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011111101100)
) lut_34_31 (
    .O(x34_y31),
    .I0(x31_y28),
    .I1(x32_y34),
    .I2(x32_y27),
    .I3(x32_y34)
);

(* keep, dont_touch *)
(* LOC = "X35/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101000100100)
) lut_35_31 (
    .O(x35_y31),
    .I0(x33_y31),
    .I1(x33_y35),
    .I2(1'b0),
    .I3(x32_y31)
);

(* keep, dont_touch *)
(* LOC = "X36/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110000000111)
) lut_36_31 (
    .O(x36_y31),
    .I0(x33_y26),
    .I1(1'b0),
    .I2(x33_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X37/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100001010110)
) lut_37_31 (
    .O(x37_y31),
    .I0(x35_y35),
    .I1(x35_y29),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X38/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100000000000)
) lut_38_31 (
    .O(x38_y31),
    .I0(x35_y36),
    .I1(x35_y36),
    .I2(x36_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X39/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100110110011)
) lut_39_31 (
    .O(x39_y31),
    .I0(1'b0),
    .I1(x37_y31),
    .I2(x37_y35),
    .I3(x37_y36)
);

(* keep, dont_touch *)
(* LOC = "X40/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100111100110)
) lut_40_31 (
    .O(x40_y31),
    .I0(x38_y33),
    .I1(x38_y30),
    .I2(x37_y26),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X41/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100100011100)
) lut_41_31 (
    .O(x41_y31),
    .I0(x38_y28),
    .I1(x38_y30),
    .I2(1'b0),
    .I3(x38_y27)
);

(* keep, dont_touch *)
(* LOC = "X42/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001111000101)
) lut_42_31 (
    .O(x42_y31),
    .I0(x39_y33),
    .I1(1'b0),
    .I2(x40_y36),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X43/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010001100011)
) lut_43_31 (
    .O(x43_y31),
    .I0(x41_y31),
    .I1(x40_y33),
    .I2(x40_y34),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X44/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110101000110)
) lut_44_31 (
    .O(x44_y31),
    .I0(x42_y29),
    .I1(x41_y34),
    .I2(x41_y29),
    .I3(x42_y26)
);

(* keep, dont_touch *)
(* LOC = "X45/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111100010000)
) lut_45_31 (
    .O(x45_y31),
    .I0(1'b0),
    .I1(x42_y27),
    .I2(x43_y26),
    .I3(x43_y26)
);

(* keep, dont_touch *)
(* LOC = "X46/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001001001110)
) lut_46_31 (
    .O(x46_y31),
    .I0(x43_y29),
    .I1(x43_y30),
    .I2(x43_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X47/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100101010001)
) lut_47_31 (
    .O(x47_y31),
    .I0(x45_y34),
    .I1(x45_y32),
    .I2(1'b0),
    .I3(x44_y31)
);

(* keep, dont_touch *)
(* LOC = "X48/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101101000001)
) lut_48_31 (
    .O(x48_y31),
    .I0(1'b0),
    .I1(x46_y34),
    .I2(1'b0),
    .I3(x46_y26)
);

(* keep, dont_touch *)
(* LOC = "X49/Y31" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101111100010)
) lut_49_31 (
    .O(x49_y31),
    .I0(x47_y32),
    .I1(x46_y26),
    .I2(x46_y34),
    .I3(x46_y32)
);

(* keep, dont_touch *)
(* LOC = "X0/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001010010000)
) lut_0_32 (
    .O(x0_y32),
    .I0(in2),
    .I1(in5),
    .I2(in9),
    .I3(in7)
);

(* keep, dont_touch *)
(* LOC = "X1/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001101001000)
) lut_1_32 (
    .O(x1_y32),
    .I0(1'b0),
    .I1(1'b0),
    .I2(in5),
    .I3(in2)
);

(* keep, dont_touch *)
(* LOC = "X2/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001000100000)
) lut_2_32 (
    .O(x2_y32),
    .I0(in0),
    .I1(in4),
    .I2(in3),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X3/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011011010011)
) lut_3_32 (
    .O(x3_y32),
    .I0(in7),
    .I1(in2),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X4/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111101000100)
) lut_4_32 (
    .O(x4_y32),
    .I0(x1_y37),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x1_y33)
);

(* keep, dont_touch *)
(* LOC = "X5/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100110110110)
) lut_5_32 (
    .O(x5_y32),
    .I0(1'b0),
    .I1(x3_y28),
    .I2(x3_y34),
    .I3(x2_y32)
);

(* keep, dont_touch *)
(* LOC = "X6/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101110000000)
) lut_6_32 (
    .O(x6_y32),
    .I0(x3_y34),
    .I1(x3_y27),
    .I2(x3_y32),
    .I3(x3_y31)
);

(* keep, dont_touch *)
(* LOC = "X7/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111101110101)
) lut_7_32 (
    .O(x7_y32),
    .I0(x5_y34),
    .I1(x4_y29),
    .I2(x4_y29),
    .I3(x4_y31)
);

(* keep, dont_touch *)
(* LOC = "X8/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010111001111)
) lut_8_32 (
    .O(x8_y32),
    .I0(x6_y35),
    .I1(x6_y29),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X9/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000000100010)
) lut_9_32 (
    .O(x9_y32),
    .I0(x7_y32),
    .I1(x6_y35),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X10/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111100010001)
) lut_10_32 (
    .O(x10_y32),
    .I0(x7_y31),
    .I1(1'b0),
    .I2(x7_y34),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X11/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100101101101)
) lut_11_32 (
    .O(x11_y32),
    .I0(x8_y29),
    .I1(x9_y37),
    .I2(x9_y35),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X12/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100101101101)
) lut_12_32 (
    .O(x12_y32),
    .I0(x9_y29),
    .I1(x10_y34),
    .I2(x10_y27),
    .I3(x10_y29)
);

(* keep, dont_touch *)
(* LOC = "X13/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101111000010)
) lut_13_32 (
    .O(x13_y32),
    .I0(1'b0),
    .I1(x11_y27),
    .I2(x11_y28),
    .I3(x11_y29)
);

(* keep, dont_touch *)
(* LOC = "X14/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000100010000)
) lut_14_32 (
    .O(x14_y32),
    .I0(x12_y35),
    .I1(x11_y34),
    .I2(x12_y27),
    .I3(x11_y28)
);

(* keep, dont_touch *)
(* LOC = "X15/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011110101110)
) lut_15_32 (
    .O(x15_y32),
    .I0(x12_y37),
    .I1(x13_y33),
    .I2(x13_y33),
    .I3(x12_y31)
);

(* keep, dont_touch *)
(* LOC = "X16/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101010110100)
) lut_16_32 (
    .O(x16_y32),
    .I0(x13_y33),
    .I1(x13_y35),
    .I2(x14_y30),
    .I3(x14_y37)
);

(* keep, dont_touch *)
(* LOC = "X17/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000001100000)
) lut_17_32 (
    .O(x17_y32),
    .I0(x14_y29),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X18/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110100011000)
) lut_18_32 (
    .O(x18_y32),
    .I0(1'b0),
    .I1(x15_y27),
    .I2(x15_y36),
    .I3(x15_y28)
);

(* keep, dont_touch *)
(* LOC = "X19/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011110011010)
) lut_19_32 (
    .O(x19_y32),
    .I0(x16_y29),
    .I1(x16_y31),
    .I2(x17_y34),
    .I3(x16_y35)
);

(* keep, dont_touch *)
(* LOC = "X20/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110110111101)
) lut_20_32 (
    .O(x20_y32),
    .I0(x17_y35),
    .I1(1'b0),
    .I2(x17_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X21/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011010000101)
) lut_21_32 (
    .O(x21_y32),
    .I0(x18_y36),
    .I1(1'b0),
    .I2(x19_y32),
    .I3(x19_y37)
);

(* keep, dont_touch *)
(* LOC = "X22/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111110001111)
) lut_22_32 (
    .O(x22_y32),
    .I0(x19_y33),
    .I1(1'b0),
    .I2(x20_y28),
    .I3(x20_y36)
);

(* keep, dont_touch *)
(* LOC = "X23/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110101101000)
) lut_23_32 (
    .O(x23_y32),
    .I0(x21_y32),
    .I1(x21_y36),
    .I2(x20_y29),
    .I3(x20_y34)
);

(* keep, dont_touch *)
(* LOC = "X24/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011110100101)
) lut_24_32 (
    .O(x24_y32),
    .I0(x21_y36),
    .I1(x21_y30),
    .I2(x21_y29),
    .I3(x21_y31)
);

(* keep, dont_touch *)
(* LOC = "X25/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000000000011)
) lut_25_32 (
    .O(x25_y32),
    .I0(x22_y27),
    .I1(1'b0),
    .I2(x22_y35),
    .I3(x23_y33)
);

(* keep, dont_touch *)
(* LOC = "X26/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101001001111)
) lut_26_32 (
    .O(x26_y32),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x24_y27),
    .I3(x23_y32)
);

(* keep, dont_touch *)
(* LOC = "X27/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111111011000)
) lut_27_32 (
    .O(x27_y32),
    .I0(x25_y35),
    .I1(x25_y30),
    .I2(x24_y34),
    .I3(x24_y28)
);

(* keep, dont_touch *)
(* LOC = "X28/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110100000110)
) lut_28_32 (
    .O(x28_y32),
    .I0(1'b0),
    .I1(x26_y28),
    .I2(x26_y27),
    .I3(x26_y27)
);

(* keep, dont_touch *)
(* LOC = "X29/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000100001011)
) lut_29_32 (
    .O(x29_y32),
    .I0(x26_y29),
    .I1(x26_y37),
    .I2(x27_y30),
    .I3(x27_y34)
);

(* keep, dont_touch *)
(* LOC = "X30/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001000101100)
) lut_30_32 (
    .O(x30_y32),
    .I0(1'b0),
    .I1(x27_y32),
    .I2(1'b0),
    .I3(x28_y33)
);

(* keep, dont_touch *)
(* LOC = "X31/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101110101000)
) lut_31_32 (
    .O(x31_y32),
    .I0(x28_y28),
    .I1(x28_y27),
    .I2(x29_y35),
    .I3(x29_y37)
);

(* keep, dont_touch *)
(* LOC = "X32/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111010001001)
) lut_32_32 (
    .O(x32_y32),
    .I0(1'b0),
    .I1(x30_y27),
    .I2(x30_y35),
    .I3(x30_y35)
);

(* keep, dont_touch *)
(* LOC = "X33/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010000000101)
) lut_33_32 (
    .O(x33_y32),
    .I0(1'b0),
    .I1(x30_y30),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X34/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011111001101)
) lut_34_32 (
    .O(x34_y32),
    .I0(x31_y35),
    .I1(1'b0),
    .I2(x31_y28),
    .I3(x31_y28)
);

(* keep, dont_touch *)
(* LOC = "X35/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011101100110)
) lut_35_32 (
    .O(x35_y32),
    .I0(x33_y30),
    .I1(x32_y28),
    .I2(x32_y33),
    .I3(x32_y29)
);

(* keep, dont_touch *)
(* LOC = "X36/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101101000010)
) lut_36_32 (
    .O(x36_y32),
    .I0(x33_y32),
    .I1(x33_y30),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X37/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100000101000)
) lut_37_32 (
    .O(x37_y32),
    .I0(1'b0),
    .I1(x34_y32),
    .I2(x34_y27),
    .I3(x35_y27)
);

(* keep, dont_touch *)
(* LOC = "X38/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010010011010)
) lut_38_32 (
    .O(x38_y32),
    .I0(x35_y37),
    .I1(1'b0),
    .I2(x35_y29),
    .I3(x35_y33)
);

(* keep, dont_touch *)
(* LOC = "X39/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011111000100)
) lut_39_32 (
    .O(x39_y32),
    .I0(x37_y27),
    .I1(x37_y31),
    .I2(x36_y37),
    .I3(x36_y27)
);

(* keep, dont_touch *)
(* LOC = "X40/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011000000101)
) lut_40_32 (
    .O(x40_y32),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x38_y29),
    .I3(x38_y35)
);

(* keep, dont_touch *)
(* LOC = "X41/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110010111001)
) lut_41_32 (
    .O(x41_y32),
    .I0(x39_y37),
    .I1(1'b0),
    .I2(x39_y32),
    .I3(x39_y29)
);

(* keep, dont_touch *)
(* LOC = "X42/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001111101001)
) lut_42_32 (
    .O(x42_y32),
    .I0(1'b0),
    .I1(x39_y30),
    .I2(x40_y32),
    .I3(x40_y36)
);

(* keep, dont_touch *)
(* LOC = "X43/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010101101111)
) lut_43_32 (
    .O(x43_y32),
    .I0(x41_y36),
    .I1(x41_y30),
    .I2(x40_y33),
    .I3(x40_y35)
);

(* keep, dont_touch *)
(* LOC = "X44/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100011110001)
) lut_44_32 (
    .O(x44_y32),
    .I0(1'b0),
    .I1(x42_y32),
    .I2(x41_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X45/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101100011011)
) lut_45_32 (
    .O(x45_y32),
    .I0(1'b0),
    .I1(x42_y36),
    .I2(1'b0),
    .I3(x43_y29)
);

(* keep, dont_touch *)
(* LOC = "X46/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111100011111)
) lut_46_32 (
    .O(x46_y32),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X47/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101110001110)
) lut_47_32 (
    .O(x47_y32),
    .I0(1'b0),
    .I1(x44_y37),
    .I2(x44_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X48/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011010100010)
) lut_48_32 (
    .O(x48_y32),
    .I0(x45_y34),
    .I1(x45_y32),
    .I2(x46_y28),
    .I3(x45_y30)
);

(* keep, dont_touch *)
(* LOC = "X49/Y32" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011010010101)
) lut_49_32 (
    .O(x49_y32),
    .I0(x46_y35),
    .I1(1'b0),
    .I2(x46_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X0/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111101000001)
) lut_0_33 (
    .O(x0_y33),
    .I0(in0),
    .I1(in2),
    .I2(in8),
    .I3(in7)
);

(* keep, dont_touch *)
(* LOC = "X1/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110110001110)
) lut_1_33 (
    .O(x1_y33),
    .I0(in8),
    .I1(in6),
    .I2(in6),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X2/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111010101110)
) lut_2_33 (
    .O(x2_y33),
    .I0(1'b0),
    .I1(1'b0),
    .I2(in9),
    .I3(in8)
);

(* keep, dont_touch *)
(* LOC = "X3/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010011000111)
) lut_3_33 (
    .O(x3_y33),
    .I0(in9),
    .I1(1'b0),
    .I2(x1_y36),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X4/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111001010100)
) lut_4_33 (
    .O(x4_y33),
    .I0(x2_y37),
    .I1(x1_y30),
    .I2(x1_y29),
    .I3(x2_y34)
);

(* keep, dont_touch *)
(* LOC = "X5/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011011111010)
) lut_5_33 (
    .O(x5_y33),
    .I0(1'b0),
    .I1(x3_y37),
    .I2(1'b0),
    .I3(x2_y31)
);

(* keep, dont_touch *)
(* LOC = "X6/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011111101101)
) lut_6_33 (
    .O(x6_y33),
    .I0(x4_y28),
    .I1(1'b0),
    .I2(x4_y28),
    .I3(x3_y31)
);

(* keep, dont_touch *)
(* LOC = "X7/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100010000000)
) lut_7_33 (
    .O(x7_y33),
    .I0(1'b0),
    .I1(x5_y29),
    .I2(x5_y36),
    .I3(x5_y32)
);

(* keep, dont_touch *)
(* LOC = "X8/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000001010100)
) lut_8_33 (
    .O(x8_y33),
    .I0(x5_y30),
    .I1(x6_y28),
    .I2(x5_y33),
    .I3(x6_y35)
);

(* keep, dont_touch *)
(* LOC = "X9/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110101101101)
) lut_9_33 (
    .O(x9_y33),
    .I0(x6_y35),
    .I1(x7_y29),
    .I2(x5_y33),
    .I3(x6_y35)
);

(* keep, dont_touch *)
(* LOC = "X10/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000100111010)
) lut_10_33 (
    .O(x10_y33),
    .I0(1'b0),
    .I1(x8_y35),
    .I2(x8_y33),
    .I3(x8_y30)
);

(* keep, dont_touch *)
(* LOC = "X11/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001100010110)
) lut_11_33 (
    .O(x11_y33),
    .I0(x8_y37),
    .I1(x8_y34),
    .I2(x9_y34),
    .I3(x8_y32)
);

(* keep, dont_touch *)
(* LOC = "X12/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111110011100)
) lut_12_33 (
    .O(x12_y33),
    .I0(1'b0),
    .I1(x10_y38),
    .I2(x10_y35),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X13/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001010111000)
) lut_13_33 (
    .O(x13_y33),
    .I0(x11_y34),
    .I1(x10_y37),
    .I2(x10_y37),
    .I3(x11_y34)
);

(* keep, dont_touch *)
(* LOC = "X14/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010010101100)
) lut_14_33 (
    .O(x14_y33),
    .I0(x11_y35),
    .I1(1'b0),
    .I2(x11_y34),
    .I3(x11_y34)
);

(* keep, dont_touch *)
(* LOC = "X15/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000100011110)
) lut_15_33 (
    .O(x15_y33),
    .I0(x13_y36),
    .I1(x13_y28),
    .I2(x12_y32),
    .I3(x13_y38)
);

(* keep, dont_touch *)
(* LOC = "X16/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110100000000)
) lut_16_33 (
    .O(x16_y33),
    .I0(x14_y29),
    .I1(x14_y29),
    .I2(1'b0),
    .I3(x13_y32)
);

(* keep, dont_touch *)
(* LOC = "X17/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110000101111)
) lut_17_33 (
    .O(x17_y33),
    .I0(x15_y32),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x15_y33)
);

(* keep, dont_touch *)
(* LOC = "X18/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101110001101)
) lut_18_33 (
    .O(x18_y33),
    .I0(1'b0),
    .I1(x15_y28),
    .I2(x15_y28),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X19/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001011011111)
) lut_19_33 (
    .O(x19_y33),
    .I0(1'b0),
    .I1(x16_y36),
    .I2(x16_y31),
    .I3(x16_y37)
);

(* keep, dont_touch *)
(* LOC = "X20/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001000011110)
) lut_20_33 (
    .O(x20_y33),
    .I0(1'b0),
    .I1(x17_y36),
    .I2(1'b0),
    .I3(x18_y34)
);

(* keep, dont_touch *)
(* LOC = "X21/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010110111110)
) lut_21_33 (
    .O(x21_y33),
    .I0(1'b0),
    .I1(x18_y38),
    .I2(x19_y37),
    .I3(x18_y32)
);

(* keep, dont_touch *)
(* LOC = "X22/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010100100100)
) lut_22_33 (
    .O(x22_y33),
    .I0(1'b0),
    .I1(x19_y37),
    .I2(1'b0),
    .I3(x20_y35)
);

(* keep, dont_touch *)
(* LOC = "X23/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001101111110)
) lut_23_33 (
    .O(x23_y33),
    .I0(x21_y29),
    .I1(1'b0),
    .I2(x20_y38),
    .I3(x20_y29)
);

(* keep, dont_touch *)
(* LOC = "X24/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100101100011)
) lut_24_33 (
    .O(x24_y33),
    .I0(1'b0),
    .I1(x21_y29),
    .I2(x21_y33),
    .I3(x21_y36)
);

(* keep, dont_touch *)
(* LOC = "X25/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100011100111)
) lut_25_33 (
    .O(x25_y33),
    .I0(1'b0),
    .I1(x22_y31),
    .I2(x22_y30),
    .I3(x23_y36)
);

(* keep, dont_touch *)
(* LOC = "X26/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000111101000)
) lut_26_33 (
    .O(x26_y33),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x23_y35),
    .I3(x23_y29)
);

(* keep, dont_touch *)
(* LOC = "X27/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101010011000)
) lut_27_33 (
    .O(x27_y33),
    .I0(x24_y32),
    .I1(x25_y29),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X28/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011100101110)
) lut_28_33 (
    .O(x28_y33),
    .I0(x25_y28),
    .I1(x26_y38),
    .I2(1'b0),
    .I3(x26_y34)
);

(* keep, dont_touch *)
(* LOC = "X29/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010011011000)
) lut_29_33 (
    .O(x29_y33),
    .I0(x26_y31),
    .I1(x27_y29),
    .I2(x27_y37),
    .I3(x27_y30)
);

(* keep, dont_touch *)
(* LOC = "X30/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010100101101)
) lut_30_33 (
    .O(x30_y33),
    .I0(x27_y29),
    .I1(x27_y28),
    .I2(x27_y31),
    .I3(x28_y33)
);

(* keep, dont_touch *)
(* LOC = "X31/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010010110110)
) lut_31_33 (
    .O(x31_y33),
    .I0(x29_y31),
    .I1(x29_y30),
    .I2(1'b0),
    .I3(x29_y37)
);

(* keep, dont_touch *)
(* LOC = "X32/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000110100001)
) lut_32_33 (
    .O(x32_y33),
    .I0(x29_y35),
    .I1(x30_y35),
    .I2(x29_y30),
    .I3(x30_y34)
);

(* keep, dont_touch *)
(* LOC = "X33/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001100111011)
) lut_33_33 (
    .O(x33_y33),
    .I0(x31_y30),
    .I1(x30_y35),
    .I2(1'b0),
    .I3(x31_y36)
);

(* keep, dont_touch *)
(* LOC = "X34/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000101010001)
) lut_34_33 (
    .O(x34_y33),
    .I0(x31_y35),
    .I1(1'b0),
    .I2(x32_y33),
    .I3(x31_y28)
);

(* keep, dont_touch *)
(* LOC = "X35/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110001100110)
) lut_35_33 (
    .O(x35_y33),
    .I0(x33_y36),
    .I1(x33_y32),
    .I2(x33_y32),
    .I3(x33_y37)
);

(* keep, dont_touch *)
(* LOC = "X36/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100110011100)
) lut_36_33 (
    .O(x36_y33),
    .I0(x33_y30),
    .I1(x34_y31),
    .I2(1'b0),
    .I3(x34_y33)
);

(* keep, dont_touch *)
(* LOC = "X37/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101000100011111)
) lut_37_33 (
    .O(x37_y33),
    .I0(x35_y29),
    .I1(1'b0),
    .I2(x34_y38),
    .I3(x34_y36)
);

(* keep, dont_touch *)
(* LOC = "X38/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100010101000)
) lut_38_33 (
    .O(x38_y33),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x36_y35),
    .I3(x35_y33)
);

(* keep, dont_touch *)
(* LOC = "X39/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100110011111)
) lut_39_33 (
    .O(x39_y33),
    .I0(1'b0),
    .I1(x36_y30),
    .I2(x36_y38),
    .I3(x36_y36)
);

(* keep, dont_touch *)
(* LOC = "X40/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100111010101)
) lut_40_33 (
    .O(x40_y33),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x37_y35),
    .I3(x38_y36)
);

(* keep, dont_touch *)
(* LOC = "X41/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101110110011)
) lut_41_33 (
    .O(x41_y33),
    .I0(x38_y33),
    .I1(1'b0),
    .I2(x39_y34),
    .I3(x38_y32)
);

(* keep, dont_touch *)
(* LOC = "X42/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011011010011)
) lut_42_33 (
    .O(x42_y33),
    .I0(x39_y30),
    .I1(x40_y38),
    .I2(1'b0),
    .I3(x39_y28)
);

(* keep, dont_touch *)
(* LOC = "X43/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111111011001)
) lut_43_33 (
    .O(x43_y33),
    .I0(x41_y29),
    .I1(1'b0),
    .I2(x41_y34),
    .I3(x40_y35)
);

(* keep, dont_touch *)
(* LOC = "X44/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000010101001)
) lut_44_33 (
    .O(x44_y33),
    .I0(1'b0),
    .I1(x42_y33),
    .I2(x41_y32),
    .I3(x42_y38)
);

(* keep, dont_touch *)
(* LOC = "X45/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010111000001)
) lut_45_33 (
    .O(x45_y33),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x42_y29),
    .I3(x43_y36)
);

(* keep, dont_touch *)
(* LOC = "X46/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111011001000)
) lut_46_33 (
    .O(x46_y33),
    .I0(x44_y38),
    .I1(x44_y33),
    .I2(x43_y32),
    .I3(x43_y33)
);

(* keep, dont_touch *)
(* LOC = "X47/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010100100010)
) lut_47_33 (
    .O(x47_y33),
    .I0(1'b0),
    .I1(x44_y30),
    .I2(x44_y29),
    .I3(x44_y33)
);

(* keep, dont_touch *)
(* LOC = "X48/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011110101010)
) lut_48_33 (
    .O(x48_y33),
    .I0(x46_y30),
    .I1(x45_y37),
    .I2(1'b0),
    .I3(x45_y36)
);

(* keep, dont_touch *)
(* LOC = "X49/Y33" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110110101011)
) lut_49_33 (
    .O(x49_y33),
    .I0(x47_y38),
    .I1(x46_y34),
    .I2(x46_y33),
    .I3(x46_y37)
);

(* keep, dont_touch *)
(* LOC = "X0/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100001100001)
) lut_0_34 (
    .O(x0_y34),
    .I0(in5),
    .I1(in0),
    .I2(in2),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X1/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010100101110)
) lut_1_34 (
    .O(x1_y34),
    .I0(in1),
    .I1(in7),
    .I2(1'b0),
    .I3(in9)
);

(* keep, dont_touch *)
(* LOC = "X2/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100010011101)
) lut_2_34 (
    .O(x2_y34),
    .I0(in1),
    .I1(in6),
    .I2(1'b0),
    .I3(in7)
);

(* keep, dont_touch *)
(* LOC = "X3/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110000001101)
) lut_3_34 (
    .O(x3_y34),
    .I0(x1_y31),
    .I1(x1_y39),
    .I2(1'b0),
    .I3(in6)
);

(* keep, dont_touch *)
(* LOC = "X4/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010111110111)
) lut_4_34 (
    .O(x4_y34),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x2_y30),
    .I3(x2_y33)
);

(* keep, dont_touch *)
(* LOC = "X5/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010110101111)
) lut_5_34 (
    .O(x5_y34),
    .I0(x3_y39),
    .I1(x3_y33),
    .I2(x3_y31),
    .I3(x2_y37)
);

(* keep, dont_touch *)
(* LOC = "X6/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101011000010)
) lut_6_34 (
    .O(x6_y34),
    .I0(x4_y33),
    .I1(x3_y37),
    .I2(x4_y34),
    .I3(x4_y39)
);

(* keep, dont_touch *)
(* LOC = "X7/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100101000011)
) lut_7_34 (
    .O(x7_y34),
    .I0(x5_y31),
    .I1(1'b0),
    .I2(x5_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X8/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111110110101)
) lut_8_34 (
    .O(x8_y34),
    .I0(x5_y32),
    .I1(x5_y34),
    .I2(1'b0),
    .I3(x5_y32)
);

(* keep, dont_touch *)
(* LOC = "X9/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010110110101)
) lut_9_34 (
    .O(x9_y34),
    .I0(x6_y39),
    .I1(x7_y35),
    .I2(1'b0),
    .I3(x5_y32)
);

(* keep, dont_touch *)
(* LOC = "X10/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011111010010)
) lut_10_34 (
    .O(x10_y34),
    .I0(x8_y33),
    .I1(x8_y33),
    .I2(1'b0),
    .I3(x8_y31)
);

(* keep, dont_touch *)
(* LOC = "X11/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001101111011)
) lut_11_34 (
    .O(x11_y34),
    .I0(x9_y38),
    .I1(x9_y33),
    .I2(x9_y37),
    .I3(x9_y29)
);

(* keep, dont_touch *)
(* LOC = "X12/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011010010100)
) lut_12_34 (
    .O(x12_y34),
    .I0(x9_y29),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x10_y35)
);

(* keep, dont_touch *)
(* LOC = "X13/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011101010011)
) lut_13_34 (
    .O(x13_y34),
    .I0(x11_y34),
    .I1(x11_y32),
    .I2(x10_y30),
    .I3(x11_y35)
);

(* keep, dont_touch *)
(* LOC = "X14/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101011001100)
) lut_14_34 (
    .O(x14_y34),
    .I0(x11_y29),
    .I1(x12_y32),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X15/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010000111110)
) lut_15_34 (
    .O(x15_y34),
    .I0(x12_y31),
    .I1(x13_y31),
    .I2(x13_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X16/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001101001101)
) lut_16_34 (
    .O(x16_y34),
    .I0(x14_y34),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x14_y30)
);

(* keep, dont_touch *)
(* LOC = "X17/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110111000000)
) lut_17_34 (
    .O(x17_y34),
    .I0(x15_y30),
    .I1(x15_y38),
    .I2(x14_y33),
    .I3(x15_y36)
);

(* keep, dont_touch *)
(* LOC = "X18/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100101010100)
) lut_18_34 (
    .O(x18_y34),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x16_y34),
    .I3(x16_y29)
);

(* keep, dont_touch *)
(* LOC = "X19/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100100011111)
) lut_19_34 (
    .O(x19_y34),
    .I0(x16_y35),
    .I1(1'b0),
    .I2(x17_y35),
    .I3(x17_y37)
);

(* keep, dont_touch *)
(* LOC = "X20/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111000100001)
) lut_20_34 (
    .O(x20_y34),
    .I0(x18_y38),
    .I1(x18_y34),
    .I2(x18_y29),
    .I3(x17_y38)
);

(* keep, dont_touch *)
(* LOC = "X21/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000111111100)
) lut_21_34 (
    .O(x21_y34),
    .I0(1'b0),
    .I1(x18_y30),
    .I2(x18_y37),
    .I3(x18_y30)
);

(* keep, dont_touch *)
(* LOC = "X22/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000100010111)
) lut_22_34 (
    .O(x22_y34),
    .I0(1'b0),
    .I1(x20_y33),
    .I2(x20_y37),
    .I3(x20_y36)
);

(* keep, dont_touch *)
(* LOC = "X23/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100011100001)
) lut_23_34 (
    .O(x23_y34),
    .I0(x21_y33),
    .I1(x20_y30),
    .I2(x21_y39),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X24/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010100011011)
) lut_24_34 (
    .O(x24_y34),
    .I0(x22_y37),
    .I1(x22_y33),
    .I2(x22_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X25/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000101110000)
) lut_25_34 (
    .O(x25_y34),
    .I0(1'b0),
    .I1(x23_y32),
    .I2(x22_y37),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X26/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110111010000)
) lut_26_34 (
    .O(x26_y34),
    .I0(1'b0),
    .I1(x24_y37),
    .I2(x24_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X27/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101000011011)
) lut_27_34 (
    .O(x27_y34),
    .I0(x25_y32),
    .I1(1'b0),
    .I2(x24_y34),
    .I3(x25_y29)
);

(* keep, dont_touch *)
(* LOC = "X28/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101000001000)
) lut_28_34 (
    .O(x28_y34),
    .I0(1'b0),
    .I1(x26_y36),
    .I2(x26_y35),
    .I3(x26_y34)
);

(* keep, dont_touch *)
(* LOC = "X29/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000110001111)
) lut_29_34 (
    .O(x29_y34),
    .I0(x26_y30),
    .I1(x27_y33),
    .I2(x26_y32),
    .I3(x26_y36)
);

(* keep, dont_touch *)
(* LOC = "X30/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111110111010)
) lut_30_34 (
    .O(x30_y34),
    .I0(x27_y36),
    .I1(x28_y36),
    .I2(x28_y31),
    .I3(x28_y38)
);

(* keep, dont_touch *)
(* LOC = "X31/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110010011100)
) lut_31_34 (
    .O(x31_y34),
    .I0(x29_y32),
    .I1(x29_y38),
    .I2(x29_y32),
    .I3(x29_y30)
);

(* keep, dont_touch *)
(* LOC = "X32/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100011100011)
) lut_32_34 (
    .O(x32_y34),
    .I0(x29_y37),
    .I1(x30_y29),
    .I2(x29_y33),
    .I3(x30_y37)
);

(* keep, dont_touch *)
(* LOC = "X33/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001111110000)
) lut_33_34 (
    .O(x33_y34),
    .I0(x30_y37),
    .I1(x31_y37),
    .I2(x31_y35),
    .I3(x31_y34)
);

(* keep, dont_touch *)
(* LOC = "X34/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100110001001)
) lut_34_34 (
    .O(x34_y34),
    .I0(x32_y32),
    .I1(x31_y30),
    .I2(1'b0),
    .I3(x31_y29)
);

(* keep, dont_touch *)
(* LOC = "X35/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100000110110)
) lut_35_34 (
    .O(x35_y34),
    .I0(x32_y39),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x32_y32)
);

(* keep, dont_touch *)
(* LOC = "X36/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011011100000)
) lut_36_34 (
    .O(x36_y34),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x33_y33),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X37/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000110100000)
) lut_37_34 (
    .O(x37_y34),
    .I0(x34_y33),
    .I1(x34_y35),
    .I2(x34_y34),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X38/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100001101010)
) lut_38_34 (
    .O(x38_y34),
    .I0(x35_y36),
    .I1(1'b0),
    .I2(x35_y38),
    .I3(x36_y37)
);

(* keep, dont_touch *)
(* LOC = "X39/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000101011110)
) lut_39_34 (
    .O(x39_y34),
    .I0(x37_y29),
    .I1(x37_y33),
    .I2(x37_y30),
    .I3(x37_y38)
);

(* keep, dont_touch *)
(* LOC = "X40/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000000110101)
) lut_40_34 (
    .O(x40_y34),
    .I0(x37_y39),
    .I1(x37_y32),
    .I2(x38_y37),
    .I3(x37_y34)
);

(* keep, dont_touch *)
(* LOC = "X41/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111011101111)
) lut_41_34 (
    .O(x41_y34),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x39_y37),
    .I3(x38_y33)
);

(* keep, dont_touch *)
(* LOC = "X42/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011111001010)
) lut_42_34 (
    .O(x42_y34),
    .I0(x40_y35),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x40_y36)
);

(* keep, dont_touch *)
(* LOC = "X43/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100001100001)
) lut_43_34 (
    .O(x43_y34),
    .I0(x40_y37),
    .I1(x40_y37),
    .I2(x41_y38),
    .I3(x41_y38)
);

(* keep, dont_touch *)
(* LOC = "X44/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100000110011)
) lut_44_34 (
    .O(x44_y34),
    .I0(x42_y32),
    .I1(x42_y29),
    .I2(x41_y37),
    .I3(x41_y33)
);

(* keep, dont_touch *)
(* LOC = "X45/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001010000100)
) lut_45_34 (
    .O(x45_y34),
    .I0(x42_y31),
    .I1(1'b0),
    .I2(x42_y30),
    .I3(x43_y34)
);

(* keep, dont_touch *)
(* LOC = "X46/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011100011111)
) lut_46_34 (
    .O(x46_y34),
    .I0(x43_y39),
    .I1(x43_y35),
    .I2(x44_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X47/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011111110001)
) lut_47_34 (
    .O(x47_y34),
    .I0(x45_y32),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x44_y39)
);

(* keep, dont_touch *)
(* LOC = "X48/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100000001010)
) lut_48_34 (
    .O(x48_y34),
    .I0(x45_y35),
    .I1(x46_y29),
    .I2(x45_y39),
    .I3(x46_y34)
);

(* keep, dont_touch *)
(* LOC = "X49/Y34" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110101111001)
) lut_49_34 (
    .O(x49_y34),
    .I0(1'b0),
    .I1(x47_y38),
    .I2(x47_y29),
    .I3(x46_y35)
);

(* keep, dont_touch *)
(* LOC = "X0/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011110010001)
) lut_0_35 (
    .O(x0_y35),
    .I0(in0),
    .I1(1'b0),
    .I2(in1),
    .I3(in1)
);

(* keep, dont_touch *)
(* LOC = "X1/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110101111111)
) lut_1_35 (
    .O(x1_y35),
    .I0(1'b0),
    .I1(in1),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X2/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111011010011)
) lut_2_35 (
    .O(x2_y35),
    .I0(in8),
    .I1(in4),
    .I2(in0),
    .I3(in5)
);

(* keep, dont_touch *)
(* LOC = "X3/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011110101110)
) lut_3_35 (
    .O(x3_y35),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x1_y39),
    .I3(in0)
);

(* keep, dont_touch *)
(* LOC = "X4/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101111111011)
) lut_4_35 (
    .O(x4_y35),
    .I0(x2_y39),
    .I1(x2_y34),
    .I2(x1_y35),
    .I3(x2_y33)
);

(* keep, dont_touch *)
(* LOC = "X5/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010000110110)
) lut_5_35 (
    .O(x5_y35),
    .I0(x3_y39),
    .I1(x2_y37),
    .I2(x2_y35),
    .I3(x2_y33)
);

(* keep, dont_touch *)
(* LOC = "X6/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000110101101)
) lut_6_35 (
    .O(x6_y35),
    .I0(x4_y40),
    .I1(x3_y34),
    .I2(1'b0),
    .I3(x3_y30)
);

(* keep, dont_touch *)
(* LOC = "X7/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011010001010)
) lut_7_35 (
    .O(x7_y35),
    .I0(x4_y36),
    .I1(x5_y30),
    .I2(1'b0),
    .I3(x5_y36)
);

(* keep, dont_touch *)
(* LOC = "X8/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010100011111)
) lut_8_35 (
    .O(x8_y35),
    .I0(x6_y30),
    .I1(x5_y37),
    .I2(x5_y40),
    .I3(x6_y37)
);

(* keep, dont_touch *)
(* LOC = "X9/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110000011001)
) lut_9_35 (
    .O(x9_y35),
    .I0(x6_y40),
    .I1(1'b0),
    .I2(x5_y40),
    .I3(x6_y37)
);

(* keep, dont_touch *)
(* LOC = "X10/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011100000001)
) lut_10_35 (
    .O(x10_y35),
    .I0(x7_y35),
    .I1(x7_y30),
    .I2(x7_y39),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X11/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000000001001)
) lut_11_35 (
    .O(x11_y35),
    .I0(x9_y36),
    .I1(x8_y34),
    .I2(x8_y30),
    .I3(x8_y31)
);

(* keep, dont_touch *)
(* LOC = "X12/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001101101010)
) lut_12_35 (
    .O(x12_y35),
    .I0(x10_y36),
    .I1(x10_y39),
    .I2(1'b0),
    .I3(x9_y35)
);

(* keep, dont_touch *)
(* LOC = "X13/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000111011000)
) lut_13_35 (
    .O(x13_y35),
    .I0(x11_y35),
    .I1(x10_y31),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X14/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010000111010)
) lut_14_35 (
    .O(x14_y35),
    .I0(x12_y33),
    .I1(x11_y40),
    .I2(x12_y32),
    .I3(x12_y35)
);

(* keep, dont_touch *)
(* LOC = "X15/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110001100000)
) lut_15_35 (
    .O(x15_y35),
    .I0(1'b0),
    .I1(x13_y36),
    .I2(x13_y38),
    .I3(x12_y36)
);

(* keep, dont_touch *)
(* LOC = "X16/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000111101110)
) lut_16_35 (
    .O(x16_y35),
    .I0(x13_y36),
    .I1(x14_y32),
    .I2(x13_y34),
    .I3(x13_y31)
);

(* keep, dont_touch *)
(* LOC = "X17/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010010111111)
) lut_17_35 (
    .O(x17_y35),
    .I0(x14_y37),
    .I1(x15_y31),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X18/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000110011101)
) lut_18_35 (
    .O(x18_y35),
    .I0(x15_y30),
    .I1(1'b0),
    .I2(x16_y34),
    .I3(x16_y33)
);

(* keep, dont_touch *)
(* LOC = "X19/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101011000111)
) lut_19_35 (
    .O(x19_y35),
    .I0(1'b0),
    .I1(x17_y30),
    .I2(1'b0),
    .I3(x17_y30)
);

(* keep, dont_touch *)
(* LOC = "X20/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111100100101)
) lut_20_35 (
    .O(x20_y35),
    .I0(x18_y38),
    .I1(x17_y37),
    .I2(x17_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X21/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111001101011)
) lut_21_35 (
    .O(x21_y35),
    .I0(x18_y31),
    .I1(x18_y40),
    .I2(x19_y39),
    .I3(x19_y40)
);

(* keep, dont_touch *)
(* LOC = "X22/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110100111000)
) lut_22_35 (
    .O(x22_y35),
    .I0(x20_y33),
    .I1(x19_y35),
    .I2(x19_y38),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X23/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111010110100)
) lut_23_35 (
    .O(x23_y35),
    .I0(x21_y39),
    .I1(x21_y32),
    .I2(x20_y39),
    .I3(x20_y31)
);

(* keep, dont_touch *)
(* LOC = "X24/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101010000111)
) lut_24_35 (
    .O(x24_y35),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x22_y33),
    .I3(x22_y32)
);

(* keep, dont_touch *)
(* LOC = "X25/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101010011011)
) lut_25_35 (
    .O(x25_y35),
    .I0(x22_y34),
    .I1(x23_y37),
    .I2(x23_y38),
    .I3(x22_y33)
);

(* keep, dont_touch *)
(* LOC = "X26/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110100100010)
) lut_26_35 (
    .O(x26_y35),
    .I0(x23_y32),
    .I1(x24_y40),
    .I2(1'b0),
    .I3(x23_y34)
);

(* keep, dont_touch *)
(* LOC = "X27/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101011111101)
) lut_27_35 (
    .O(x27_y35),
    .I0(x25_y37),
    .I1(x24_y31),
    .I2(x25_y35),
    .I3(x24_y35)
);

(* keep, dont_touch *)
(* LOC = "X28/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100001011000)
) lut_28_35 (
    .O(x28_y35),
    .I0(x26_y34),
    .I1(x26_y39),
    .I2(x25_y34),
    .I3(x25_y30)
);

(* keep, dont_touch *)
(* LOC = "X29/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011000111001)
) lut_29_35 (
    .O(x29_y35),
    .I0(1'b0),
    .I1(x27_y33),
    .I2(x27_y35),
    .I3(x26_y40)
);

(* keep, dont_touch *)
(* LOC = "X30/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000010010101)
) lut_30_35 (
    .O(x30_y35),
    .I0(x28_y35),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x28_y30)
);

(* keep, dont_touch *)
(* LOC = "X31/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111011011011)
) lut_31_35 (
    .O(x31_y35),
    .I0(x29_y37),
    .I1(x28_y31),
    .I2(x28_y39),
    .I3(x29_y35)
);

(* keep, dont_touch *)
(* LOC = "X32/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000110110101)
) lut_32_35 (
    .O(x32_y35),
    .I0(x30_y37),
    .I1(x29_y36),
    .I2(x30_y30),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X33/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010010010000)
) lut_33_35 (
    .O(x33_y35),
    .I0(1'b0),
    .I1(x31_y33),
    .I2(x31_y37),
    .I3(x31_y32)
);

(* keep, dont_touch *)
(* LOC = "X34/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111100011101)
) lut_34_35 (
    .O(x34_y35),
    .I0(x31_y39),
    .I1(x31_y31),
    .I2(x31_y32),
    .I3(x31_y34)
);

(* keep, dont_touch *)
(* LOC = "X35/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110101110110)
) lut_35_35 (
    .O(x35_y35),
    .I0(x32_y32),
    .I1(x33_y38),
    .I2(1'b0),
    .I3(x33_y34)
);

(* keep, dont_touch *)
(* LOC = "X36/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110000100010)
) lut_36_35 (
    .O(x36_y35),
    .I0(x33_y36),
    .I1(x34_y32),
    .I2(1'b0),
    .I3(x33_y37)
);

(* keep, dont_touch *)
(* LOC = "X37/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000100001010)
) lut_37_35 (
    .O(x37_y35),
    .I0(x35_y30),
    .I1(x34_y32),
    .I2(x35_y33),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X38/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101110000111)
) lut_38_35 (
    .O(x38_y35),
    .I0(1'b0),
    .I1(x36_y38),
    .I2(x35_y39),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X39/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101000100010)
) lut_39_35 (
    .O(x39_y35),
    .I0(x36_y38),
    .I1(1'b0),
    .I2(x37_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X40/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110111101101)
) lut_40_35 (
    .O(x40_y35),
    .I0(x38_y33),
    .I1(1'b0),
    .I2(x38_y38),
    .I3(x38_y32)
);

(* keep, dont_touch *)
(* LOC = "X41/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000110011110)
) lut_41_35 (
    .O(x41_y35),
    .I0(x38_y37),
    .I1(x39_y32),
    .I2(x39_y39),
    .I3(x38_y32)
);

(* keep, dont_touch *)
(* LOC = "X42/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101010011000)
) lut_42_35 (
    .O(x42_y35),
    .I0(x39_y31),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x39_y32)
);

(* keep, dont_touch *)
(* LOC = "X43/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101101001110)
) lut_43_35 (
    .O(x43_y35),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x40_y37)
);

(* keep, dont_touch *)
(* LOC = "X44/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011010110010)
) lut_44_35 (
    .O(x44_y35),
    .I0(x42_y32),
    .I1(x42_y39),
    .I2(x41_y33),
    .I3(x41_y38)
);

(* keep, dont_touch *)
(* LOC = "X45/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110110001111)
) lut_45_35 (
    .O(x45_y35),
    .I0(x43_y30),
    .I1(1'b0),
    .I2(x43_y40),
    .I3(x42_y34)
);

(* keep, dont_touch *)
(* LOC = "X46/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111110101010)
) lut_46_35 (
    .O(x46_y35),
    .I0(x43_y37),
    .I1(1'b0),
    .I2(x43_y34),
    .I3(x44_y34)
);

(* keep, dont_touch *)
(* LOC = "X47/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100000110100)
) lut_47_35 (
    .O(x47_y35),
    .I0(1'b0),
    .I1(x45_y31),
    .I2(x44_y39),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X48/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111111011000)
) lut_48_35 (
    .O(x48_y35),
    .I0(x46_y31),
    .I1(x45_y36),
    .I2(x45_y35),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X49/Y35" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000111110101)
) lut_49_35 (
    .O(x49_y35),
    .I0(x46_y31),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x47_y36)
);

(* keep, dont_touch *)
(* LOC = "X0/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111011000001)
) lut_0_36 (
    .O(x0_y36),
    .I0(in8),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X1/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010011100101)
) lut_1_36 (
    .O(x1_y36),
    .I0(in6),
    .I1(in8),
    .I2(1'b0),
    .I3(in6)
);

(* keep, dont_touch *)
(* LOC = "X2/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010011100001)
) lut_2_36 (
    .O(x2_y36),
    .I0(in9),
    .I1(in1),
    .I2(in1),
    .I3(in1)
);

(* keep, dont_touch *)
(* LOC = "X3/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111010001001)
) lut_3_36 (
    .O(x3_y36),
    .I0(in8),
    .I1(in4),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X4/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110000101011)
) lut_4_36 (
    .O(x4_y36),
    .I0(x1_y39),
    .I1(x1_y33),
    .I2(1'b0),
    .I3(x1_y34)
);

(* keep, dont_touch *)
(* LOC = "X5/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111000001001)
) lut_5_36 (
    .O(x5_y36),
    .I0(x2_y33),
    .I1(x2_y39),
    .I2(x2_y37),
    .I3(x2_y35)
);

(* keep, dont_touch *)
(* LOC = "X6/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100010001001)
) lut_6_36 (
    .O(x6_y36),
    .I0(x3_y40),
    .I1(x4_y36),
    .I2(x3_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X7/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001100100011)
) lut_7_36 (
    .O(x7_y36),
    .I0(x4_y36),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x4_y38)
);

(* keep, dont_touch *)
(* LOC = "X8/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110011000001)
) lut_8_36 (
    .O(x8_y36),
    .I0(1'b0),
    .I1(x5_y40),
    .I2(x5_y36),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X9/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000001001000)
) lut_9_36 (
    .O(x9_y36),
    .I0(x6_y38),
    .I1(x6_y37),
    .I2(x5_y36),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X10/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001101010110)
) lut_10_36 (
    .O(x10_y36),
    .I0(x8_y41),
    .I1(x7_y34),
    .I2(x7_y37),
    .I3(x8_y40)
);

(* keep, dont_touch *)
(* LOC = "X11/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110110110110)
) lut_11_36 (
    .O(x11_y36),
    .I0(x8_y31),
    .I1(x9_y32),
    .I2(x9_y35),
    .I3(x8_y40)
);

(* keep, dont_touch *)
(* LOC = "X12/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100100101111)
) lut_12_36 (
    .O(x12_y36),
    .I0(x9_y41),
    .I1(x9_y39),
    .I2(x9_y40),
    .I3(x10_y35)
);

(* keep, dont_touch *)
(* LOC = "X13/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001000111010)
) lut_13_36 (
    .O(x13_y36),
    .I0(x11_y31),
    .I1(x10_y35),
    .I2(x10_y33),
    .I3(x11_y41)
);

(* keep, dont_touch *)
(* LOC = "X14/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011000010010)
) lut_14_36 (
    .O(x14_y36),
    .I0(x11_y32),
    .I1(x11_y31),
    .I2(x11_y34),
    .I3(x11_y32)
);

(* keep, dont_touch *)
(* LOC = "X15/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010010011001)
) lut_15_36 (
    .O(x15_y36),
    .I0(1'b0),
    .I1(x13_y40),
    .I2(x12_y40),
    .I3(x13_y32)
);

(* keep, dont_touch *)
(* LOC = "X16/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011001100100)
) lut_16_36 (
    .O(x16_y36),
    .I0(1'b0),
    .I1(x14_y31),
    .I2(1'b0),
    .I3(x14_y33)
);

(* keep, dont_touch *)
(* LOC = "X17/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001111001011)
) lut_17_36 (
    .O(x17_y36),
    .I0(x14_y33),
    .I1(x14_y31),
    .I2(x15_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X18/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101011000110)
) lut_18_36 (
    .O(x18_y36),
    .I0(1'b0),
    .I1(x16_y32),
    .I2(1'b0),
    .I3(x16_y41)
);

(* keep, dont_touch *)
(* LOC = "X19/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100111010111)
) lut_19_36 (
    .O(x19_y36),
    .I0(1'b0),
    .I1(x17_y31),
    .I2(x16_y39),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X20/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000110111101)
) lut_20_36 (
    .O(x20_y36),
    .I0(x17_y33),
    .I1(x17_y39),
    .I2(x18_y33),
    .I3(x17_y41)
);

(* keep, dont_touch *)
(* LOC = "X21/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101101111010)
) lut_21_36 (
    .O(x21_y36),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x18_y41)
);

(* keep, dont_touch *)
(* LOC = "X22/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100100101001)
) lut_22_36 (
    .O(x22_y36),
    .I0(x20_y37),
    .I1(1'b0),
    .I2(x20_y38),
    .I3(x19_y33)
);

(* keep, dont_touch *)
(* LOC = "X23/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010111011000)
) lut_23_36 (
    .O(x23_y36),
    .I0(x20_y41),
    .I1(1'b0),
    .I2(x20_y32),
    .I3(x20_y36)
);

(* keep, dont_touch *)
(* LOC = "X24/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100000011011)
) lut_24_36 (
    .O(x24_y36),
    .I0(x22_y35),
    .I1(x21_y33),
    .I2(x22_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X25/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101001110110)
) lut_25_36 (
    .O(x25_y36),
    .I0(x23_y39),
    .I1(x23_y41),
    .I2(1'b0),
    .I3(x22_y41)
);

(* keep, dont_touch *)
(* LOC = "X26/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100010100101)
) lut_26_36 (
    .O(x26_y36),
    .I0(x24_y39),
    .I1(x23_y38),
    .I2(1'b0),
    .I3(x23_y32)
);

(* keep, dont_touch *)
(* LOC = "X27/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101100010001)
) lut_27_36 (
    .O(x27_y36),
    .I0(x24_y34),
    .I1(x24_y38),
    .I2(x25_y31),
    .I3(x25_y37)
);

(* keep, dont_touch *)
(* LOC = "X28/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100011011111)
) lut_28_36 (
    .O(x28_y36),
    .I0(x25_y39),
    .I1(1'b0),
    .I2(x26_y40),
    .I3(x25_y32)
);

(* keep, dont_touch *)
(* LOC = "X29/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010111011011)
) lut_29_36 (
    .O(x29_y36),
    .I0(x27_y36),
    .I1(x27_y32),
    .I2(x27_y31),
    .I3(x27_y36)
);

(* keep, dont_touch *)
(* LOC = "X30/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111001110111)
) lut_30_36 (
    .O(x30_y36),
    .I0(x28_y40),
    .I1(x27_y39),
    .I2(1'b0),
    .I3(x28_y34)
);

(* keep, dont_touch *)
(* LOC = "X31/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111010100110)
) lut_31_36 (
    .O(x31_y36),
    .I0(x29_y32),
    .I1(x29_y32),
    .I2(x28_y31),
    .I3(x28_y33)
);

(* keep, dont_touch *)
(* LOC = "X32/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011000100100)
) lut_32_36 (
    .O(x32_y36),
    .I0(x30_y38),
    .I1(x30_y40),
    .I2(1'b0),
    .I3(x29_y41)
);

(* keep, dont_touch *)
(* LOC = "X33/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101110110001)
) lut_33_36 (
    .O(x33_y36),
    .I0(x30_y41),
    .I1(x31_y40),
    .I2(x31_y38),
    .I3(x30_y32)
);

(* keep, dont_touch *)
(* LOC = "X34/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100110100000)
) lut_34_36 (
    .O(x34_y36),
    .I0(x32_y40),
    .I1(x32_y40),
    .I2(x32_y34),
    .I3(x32_y32)
);

(* keep, dont_touch *)
(* LOC = "X35/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101000110111)
) lut_35_36 (
    .O(x35_y36),
    .I0(x32_y33),
    .I1(x32_y31),
    .I2(x32_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X36/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110101001011)
) lut_36_36 (
    .O(x36_y36),
    .I0(x33_y35),
    .I1(x33_y32),
    .I2(x34_y35),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X37/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101010101000)
) lut_37_36 (
    .O(x37_y36),
    .I0(x34_y39),
    .I1(x35_y35),
    .I2(x35_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X38/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010011100001)
) lut_38_36 (
    .O(x38_y36),
    .I0(1'b0),
    .I1(x35_y34),
    .I2(x35_y34),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X39/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101001010100)
) lut_39_36 (
    .O(x39_y36),
    .I0(x36_y31),
    .I1(x37_y39),
    .I2(x36_y31),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X40/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101001101101)
) lut_40_36 (
    .O(x40_y36),
    .I0(x37_y31),
    .I1(x38_y35),
    .I2(x37_y41),
    .I3(x38_y40)
);

(* keep, dont_touch *)
(* LOC = "X41/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110111010101)
) lut_41_36 (
    .O(x41_y36),
    .I0(x38_y39),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x39_y31)
);

(* keep, dont_touch *)
(* LOC = "X42/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000110001101)
) lut_42_36 (
    .O(x42_y36),
    .I0(1'b0),
    .I1(x39_y35),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X43/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101100000101)
) lut_43_36 (
    .O(x43_y36),
    .I0(x40_y38),
    .I1(x40_y39),
    .I2(x40_y38),
    .I3(x41_y33)
);

(* keep, dont_touch *)
(* LOC = "X44/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101000011100)
) lut_44_36 (
    .O(x44_y36),
    .I0(1'b0),
    .I1(x42_y37),
    .I2(x42_y37),
    .I3(x42_y35)
);

(* keep, dont_touch *)
(* LOC = "X45/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111010010000)
) lut_45_36 (
    .O(x45_y36),
    .I0(x43_y40),
    .I1(1'b0),
    .I2(x43_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X46/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001001000001)
) lut_46_36 (
    .O(x46_y36),
    .I0(x43_y32),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X47/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011010010000)
) lut_47_36 (
    .O(x47_y36),
    .I0(x44_y39),
    .I1(x44_y33),
    .I2(x44_y35),
    .I3(x45_y34)
);

(* keep, dont_touch *)
(* LOC = "X48/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110010001010)
) lut_48_36 (
    .O(x48_y36),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x46_y37),
    .I3(x46_y41)
);

(* keep, dont_touch *)
(* LOC = "X49/Y36" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110011001100)
) lut_49_36 (
    .O(x49_y36),
    .I0(x46_y38),
    .I1(x47_y34),
    .I2(x47_y38),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X0/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001010011100)
) lut_0_37 (
    .O(x0_y37),
    .I0(in3),
    .I1(in4),
    .I2(1'b0),
    .I3(in2)
);

(* keep, dont_touch *)
(* LOC = "X1/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011001011111)
) lut_1_37 (
    .O(x1_y37),
    .I0(in4),
    .I1(in0),
    .I2(in5),
    .I3(in5)
);

(* keep, dont_touch *)
(* LOC = "X2/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101001110010)
) lut_2_37 (
    .O(x2_y37),
    .I0(1'b0),
    .I1(in2),
    .I2(in7),
    .I3(in2)
);

(* keep, dont_touch *)
(* LOC = "X3/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110101100100)
) lut_3_37 (
    .O(x3_y37),
    .I0(x1_y35),
    .I1(x1_y36),
    .I2(1'b0),
    .I3(in5)
);

(* keep, dont_touch *)
(* LOC = "X4/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100000000011)
) lut_4_37 (
    .O(x4_y37),
    .I0(x1_y39),
    .I1(x2_y37),
    .I2(x1_y34),
    .I3(x1_y32)
);

(* keep, dont_touch *)
(* LOC = "X5/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100110110111)
) lut_5_37 (
    .O(x5_y37),
    .I0(x2_y42),
    .I1(1'b0),
    .I2(x2_y37),
    .I3(x2_y40)
);

(* keep, dont_touch *)
(* LOC = "X6/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001101101001)
) lut_6_37 (
    .O(x6_y37),
    .I0(x3_y39),
    .I1(1'b0),
    .I2(x4_y34),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X7/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110101101100)
) lut_7_37 (
    .O(x7_y37),
    .I0(x4_y32),
    .I1(x5_y42),
    .I2(x4_y33),
    .I3(x5_y36)
);

(* keep, dont_touch *)
(* LOC = "X8/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100011111010)
) lut_8_37 (
    .O(x8_y37),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X9/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010101010001)
) lut_9_37 (
    .O(x9_y37),
    .I0(1'b0),
    .I1(x6_y40),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X10/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011111010100)
) lut_10_37 (
    .O(x10_y37),
    .I0(x8_y41),
    .I1(x7_y35),
    .I2(x7_y39),
    .I3(x7_y36)
);

(* keep, dont_touch *)
(* LOC = "X11/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101111100010)
) lut_11_37 (
    .O(x11_y37),
    .I0(1'b0),
    .I1(x8_y34),
    .I2(x8_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X12/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001101010111)
) lut_12_37 (
    .O(x12_y37),
    .I0(1'b0),
    .I1(x9_y37),
    .I2(x10_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X13/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010001101101)
) lut_13_37 (
    .O(x13_y37),
    .I0(x10_y40),
    .I1(x11_y40),
    .I2(x10_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X14/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010000011111)
) lut_14_37 (
    .O(x14_y37),
    .I0(x12_y36),
    .I1(x12_y33),
    .I2(x12_y41),
    .I3(x11_y37)
);

(* keep, dont_touch *)
(* LOC = "X15/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000000101000)
) lut_15_37 (
    .O(x15_y37),
    .I0(x12_y37),
    .I1(x12_y36),
    .I2(x12_y37),
    .I3(x12_y39)
);

(* keep, dont_touch *)
(* LOC = "X16/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110101101101)
) lut_16_37 (
    .O(x16_y37),
    .I0(x13_y37),
    .I1(x13_y41),
    .I2(x13_y33),
    .I3(x13_y40)
);

(* keep, dont_touch *)
(* LOC = "X17/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000010110010)
) lut_17_37 (
    .O(x17_y37),
    .I0(1'b0),
    .I1(x15_y34),
    .I2(x14_y41),
    .I3(x15_y38)
);

(* keep, dont_touch *)
(* LOC = "X18/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111100110011)
) lut_18_37 (
    .O(x18_y37),
    .I0(x15_y32),
    .I1(x16_y41),
    .I2(x16_y33),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X19/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100111000011)
) lut_19_37 (
    .O(x19_y37),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x17_y42),
    .I3(x17_y39)
);

(* keep, dont_touch *)
(* LOC = "X20/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110000011010)
) lut_20_37 (
    .O(x20_y37),
    .I0(x18_y32),
    .I1(x18_y38),
    .I2(x17_y41),
    .I3(x17_y41)
);

(* keep, dont_touch *)
(* LOC = "X21/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010010101001)
) lut_21_37 (
    .O(x21_y37),
    .I0(x18_y40),
    .I1(x19_y40),
    .I2(x19_y39),
    .I3(x19_y42)
);

(* keep, dont_touch *)
(* LOC = "X22/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101000111011)
) lut_22_37 (
    .O(x22_y37),
    .I0(x19_y35),
    .I1(x19_y37),
    .I2(1'b0),
    .I3(x19_y33)
);

(* keep, dont_touch *)
(* LOC = "X23/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111011101011)
) lut_23_37 (
    .O(x23_y37),
    .I0(x20_y40),
    .I1(x20_y34),
    .I2(x20_y38),
    .I3(x21_y38)
);

(* keep, dont_touch *)
(* LOC = "X24/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011111000101)
) lut_24_37 (
    .O(x24_y37),
    .I0(x22_y38),
    .I1(x21_y39),
    .I2(1'b0),
    .I3(x22_y36)
);

(* keep, dont_touch *)
(* LOC = "X25/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100000011111)
) lut_25_37 (
    .O(x25_y37),
    .I0(x23_y33),
    .I1(x23_y36),
    .I2(x23_y32),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X26/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111100100110)
) lut_26_37 (
    .O(x26_y37),
    .I0(x23_y33),
    .I1(1'b0),
    .I2(x24_y32),
    .I3(x23_y41)
);

(* keep, dont_touch *)
(* LOC = "X27/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101101110011)
) lut_27_37 (
    .O(x27_y37),
    .I0(x25_y33),
    .I1(1'b0),
    .I2(x24_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X28/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100000110011)
) lut_28_37 (
    .O(x28_y37),
    .I0(x25_y35),
    .I1(1'b0),
    .I2(x25_y36),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X29/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100101110010)
) lut_29_37 (
    .O(x29_y37),
    .I0(x26_y34),
    .I1(1'b0),
    .I2(x26_y39),
    .I3(x26_y33)
);

(* keep, dont_touch *)
(* LOC = "X30/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110101000000)
) lut_30_37 (
    .O(x30_y37),
    .I0(x28_y40),
    .I1(x28_y32),
    .I2(x27_y38),
    .I3(x27_y42)
);

(* keep, dont_touch *)
(* LOC = "X31/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111111000101)
) lut_31_37 (
    .O(x31_y37),
    .I0(1'b0),
    .I1(x28_y40),
    .I2(x29_y39),
    .I3(x29_y38)
);

(* keep, dont_touch *)
(* LOC = "X32/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000101011001)
) lut_32_37 (
    .O(x32_y37),
    .I0(x29_y36),
    .I1(x29_y41),
    .I2(x29_y38),
    .I3(x30_y40)
);

(* keep, dont_touch *)
(* LOC = "X33/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000011010100)
) lut_33_37 (
    .O(x33_y37),
    .I0(1'b0),
    .I1(x31_y35),
    .I2(x31_y41),
    .I3(x31_y42)
);

(* keep, dont_touch *)
(* LOC = "X34/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010000101001)
) lut_34_37 (
    .O(x34_y37),
    .I0(x31_y37),
    .I1(1'b0),
    .I2(x32_y40),
    .I3(x32_y33)
);

(* keep, dont_touch *)
(* LOC = "X35/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100100111110)
) lut_35_37 (
    .O(x35_y37),
    .I0(x32_y35),
    .I1(1'b0),
    .I2(x32_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X36/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110101110011)
) lut_36_37 (
    .O(x36_y37),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x34_y35),
    .I3(x34_y37)
);

(* keep, dont_touch *)
(* LOC = "X37/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101000111000)
) lut_37_37 (
    .O(x37_y37),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x35_y38),
    .I3(x34_y33)
);

(* keep, dont_touch *)
(* LOC = "X38/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101110100101)
) lut_38_37 (
    .O(x38_y37),
    .I0(1'b0),
    .I1(x36_y42),
    .I2(1'b0),
    .I3(x36_y38)
);

(* keep, dont_touch *)
(* LOC = "X39/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111101110001)
) lut_39_37 (
    .O(x39_y37),
    .I0(1'b0),
    .I1(x36_y32),
    .I2(x36_y38),
    .I3(x36_y40)
);

(* keep, dont_touch *)
(* LOC = "X40/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000101111011)
) lut_40_37 (
    .O(x40_y37),
    .I0(1'b0),
    .I1(x37_y32),
    .I2(x38_y41),
    .I3(x37_y39)
);

(* keep, dont_touch *)
(* LOC = "X41/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101010001100)
) lut_41_37 (
    .O(x41_y37),
    .I0(x39_y33),
    .I1(x38_y35),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X42/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100010101111)
) lut_42_37 (
    .O(x42_y37),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x40_y42),
    .I3(x39_y34)
);

(* keep, dont_touch *)
(* LOC = "X43/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100000100001)
) lut_43_37 (
    .O(x43_y37),
    .I0(x40_y35),
    .I1(x40_y42),
    .I2(x40_y34),
    .I3(x41_y38)
);

(* keep, dont_touch *)
(* LOC = "X44/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100110011110)
) lut_44_37 (
    .O(x44_y37),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x42_y42),
    .I3(x42_y32)
);

(* keep, dont_touch *)
(* LOC = "X45/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011000000010)
) lut_45_37 (
    .O(x45_y37),
    .I0(x43_y42),
    .I1(x42_y34),
    .I2(1'b0),
    .I3(x42_y35)
);

(* keep, dont_touch *)
(* LOC = "X46/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110011110101)
) lut_46_37 (
    .O(x46_y37),
    .I0(1'b0),
    .I1(x43_y39),
    .I2(x44_y38),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X47/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000110010000)
) lut_47_37 (
    .O(x47_y37),
    .I0(x45_y32),
    .I1(1'b0),
    .I2(x45_y35),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X48/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011100000111)
) lut_48_37 (
    .O(x48_y37),
    .I0(x46_y33),
    .I1(x45_y40),
    .I2(x45_y40),
    .I3(x46_y32)
);

(* keep, dont_touch *)
(* LOC = "X49/Y37" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101011001110)
) lut_49_37 (
    .O(x49_y37),
    .I0(x46_y32),
    .I1(x46_y33),
    .I2(x47_y38),
    .I3(x46_y37)
);

(* keep, dont_touch *)
(* LOC = "X0/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011010110011)
) lut_0_38 (
    .O(x0_y38),
    .I0(in3),
    .I1(in3),
    .I2(in7),
    .I3(in6)
);

(* keep, dont_touch *)
(* LOC = "X1/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001111011110)
) lut_1_38 (
    .O(x1_y38),
    .I0(in2),
    .I1(in9),
    .I2(1'b0),
    .I3(in8)
);

(* keep, dont_touch *)
(* LOC = "X2/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100111001110)
) lut_2_38 (
    .O(x2_y38),
    .I0(in8),
    .I1(in5),
    .I2(in3),
    .I3(in7)
);

(* keep, dont_touch *)
(* LOC = "X3/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011010011111)
) lut_3_38 (
    .O(x3_y38),
    .I0(in4),
    .I1(x1_y33),
    .I2(in7),
    .I3(in2)
);

(* keep, dont_touch *)
(* LOC = "X4/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000000111101)
) lut_4_38 (
    .O(x4_y38),
    .I0(x2_y36),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x1_y35)
);

(* keep, dont_touch *)
(* LOC = "X5/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010100100100)
) lut_5_38 (
    .O(x5_y38),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x3_y40),
    .I3(x3_y38)
);

(* keep, dont_touch *)
(* LOC = "X6/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010000110100)
) lut_6_38 (
    .O(x6_y38),
    .I0(x3_y42),
    .I1(x4_y42),
    .I2(1'b0),
    .I3(x4_y41)
);

(* keep, dont_touch *)
(* LOC = "X7/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001000011110)
) lut_7_38 (
    .O(x7_y38),
    .I0(x4_y40),
    .I1(x5_y43),
    .I2(x4_y35),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X8/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010100101010)
) lut_8_38 (
    .O(x8_y38),
    .I0(x5_y38),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x5_y38)
);

(* keep, dont_touch *)
(* LOC = "X9/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001010010110)
) lut_9_38 (
    .O(x9_y38),
    .I0(x7_y33),
    .I1(x7_y38),
    .I2(1'b0),
    .I3(x5_y38)
);

(* keep, dont_touch *)
(* LOC = "X10/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111100110000)
) lut_10_38 (
    .O(x10_y38),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x8_y38),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X11/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110000110101)
) lut_11_38 (
    .O(x11_y38),
    .I0(x8_y33),
    .I1(x8_y33),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X12/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011000110101)
) lut_12_38 (
    .O(x12_y38),
    .I0(1'b0),
    .I1(x10_y42),
    .I2(1'b0),
    .I3(x9_y35)
);

(* keep, dont_touch *)
(* LOC = "X13/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110100010000)
) lut_13_38 (
    .O(x13_y38),
    .I0(x10_y38),
    .I1(x10_y33),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X14/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001010010010)
) lut_14_38 (
    .O(x14_y38),
    .I0(1'b0),
    .I1(x11_y37),
    .I2(x12_y41),
    .I3(x11_y37)
);

(* keep, dont_touch *)
(* LOC = "X15/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101011101001)
) lut_15_38 (
    .O(x15_y38),
    .I0(1'b0),
    .I1(x13_y38),
    .I2(x12_y39),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X16/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011000100010)
) lut_16_38 (
    .O(x16_y38),
    .I0(x13_y35),
    .I1(x14_y41),
    .I2(x13_y38),
    .I3(x14_y37)
);

(* keep, dont_touch *)
(* LOC = "X17/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101100110111)
) lut_17_38 (
    .O(x17_y38),
    .I0(x14_y43),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x14_y39)
);

(* keep, dont_touch *)
(* LOC = "X18/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010100000110)
) lut_18_38 (
    .O(x18_y38),
    .I0(x15_y36),
    .I1(1'b0),
    .I2(x15_y40),
    .I3(x16_y38)
);

(* keep, dont_touch *)
(* LOC = "X19/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110000100110111)
) lut_19_38 (
    .O(x19_y38),
    .I0(1'b0),
    .I1(x16_y43),
    .I2(x17_y39),
    .I3(x17_y37)
);

(* keep, dont_touch *)
(* LOC = "X20/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011110000100)
) lut_20_38 (
    .O(x20_y38),
    .I0(x17_y37),
    .I1(1'b0),
    .I2(x17_y36),
    .I3(x17_y39)
);

(* keep, dont_touch *)
(* LOC = "X21/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110100011011)
) lut_21_38 (
    .O(x21_y38),
    .I0(x19_y43),
    .I1(x19_y38),
    .I2(x19_y33),
    .I3(x19_y42)
);

(* keep, dont_touch *)
(* LOC = "X22/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010010100100)
) lut_22_38 (
    .O(x22_y38),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x19_y35),
    .I3(x19_y41)
);

(* keep, dont_touch *)
(* LOC = "X23/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101011001001)
) lut_23_38 (
    .O(x23_y38),
    .I0(x21_y39),
    .I1(x20_y40),
    .I2(x21_y43),
    .I3(x21_y38)
);

(* keep, dont_touch *)
(* LOC = "X24/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111111100101)
) lut_24_38 (
    .O(x24_y38),
    .I0(x21_y35),
    .I1(x21_y33),
    .I2(1'b0),
    .I3(x21_y41)
);

(* keep, dont_touch *)
(* LOC = "X25/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111111100100)
) lut_25_38 (
    .O(x25_y38),
    .I0(x23_y37),
    .I1(x22_y34),
    .I2(x23_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X26/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000011110010)
) lut_26_38 (
    .O(x26_y38),
    .I0(x23_y33),
    .I1(x24_y37),
    .I2(x23_y34),
    .I3(x23_y43)
);

(* keep, dont_touch *)
(* LOC = "X27/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101000010110)
) lut_27_38 (
    .O(x27_y38),
    .I0(x24_y37),
    .I1(x25_y37),
    .I2(x25_y43),
    .I3(x24_y41)
);

(* keep, dont_touch *)
(* LOC = "X28/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010000010011)
) lut_28_38 (
    .O(x28_y38),
    .I0(1'b0),
    .I1(x25_y33),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X29/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001101110100)
) lut_29_38 (
    .O(x29_y38),
    .I0(x26_y35),
    .I1(x26_y35),
    .I2(x27_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X30/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100000000100)
) lut_30_38 (
    .O(x30_y38),
    .I0(x28_y37),
    .I1(x28_y37),
    .I2(1'b0),
    .I3(x27_y37)
);

(* keep, dont_touch *)
(* LOC = "X31/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101000000100)
) lut_31_38 (
    .O(x31_y38),
    .I0(x29_y41),
    .I1(x28_y33),
    .I2(x29_y41),
    .I3(x28_y42)
);

(* keep, dont_touch *)
(* LOC = "X32/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100010101001)
) lut_32_38 (
    .O(x32_y38),
    .I0(x29_y42),
    .I1(x29_y39),
    .I2(x30_y38),
    .I3(x30_y34)
);

(* keep, dont_touch *)
(* LOC = "X33/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010000110001)
) lut_33_38 (
    .O(x33_y38),
    .I0(x31_y41),
    .I1(1'b0),
    .I2(x30_y35),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X34/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110000100011)
) lut_34_38 (
    .O(x34_y38),
    .I0(x32_y39),
    .I1(x31_y35),
    .I2(x32_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X35/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000000111011)
) lut_35_38 (
    .O(x35_y38),
    .I0(x33_y33),
    .I1(x33_y40),
    .I2(x32_y41),
    .I3(x32_y34)
);

(* keep, dont_touch *)
(* LOC = "X36/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110100000001)
) lut_36_38 (
    .O(x36_y38),
    .I0(x33_y34),
    .I1(x33_y39),
    .I2(x34_y39),
    .I3(x33_y37)
);

(* keep, dont_touch *)
(* LOC = "X37/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011010000000)
) lut_37_38 (
    .O(x37_y38),
    .I0(x34_y39),
    .I1(1'b0),
    .I2(x34_y38),
    .I3(x35_y36)
);

(* keep, dont_touch *)
(* LOC = "X38/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100100010110)
) lut_38_38 (
    .O(x38_y38),
    .I0(x36_y39),
    .I1(x36_y35),
    .I2(x36_y42),
    .I3(x35_y40)
);

(* keep, dont_touch *)
(* LOC = "X39/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010001110100)
) lut_39_38 (
    .O(x39_y38),
    .I0(x37_y38),
    .I1(x36_y35),
    .I2(x36_y37),
    .I3(x36_y37)
);

(* keep, dont_touch *)
(* LOC = "X40/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011011100000)
) lut_40_38 (
    .O(x40_y38),
    .I0(x38_y40),
    .I1(x38_y34),
    .I2(x38_y37),
    .I3(x38_y41)
);

(* keep, dont_touch *)
(* LOC = "X41/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111000001000)
) lut_41_38 (
    .O(x41_y38),
    .I0(x39_y37),
    .I1(x38_y40),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X42/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000110000111)
) lut_42_38 (
    .O(x42_y38),
    .I0(x40_y39),
    .I1(1'b0),
    .I2(x40_y43),
    .I3(x40_y42)
);

(* keep, dont_touch *)
(* LOC = "X43/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001001111111)
) lut_43_38 (
    .O(x43_y38),
    .I0(x40_y41),
    .I1(x41_y40),
    .I2(x41_y37),
    .I3(x40_y35)
);

(* keep, dont_touch *)
(* LOC = "X44/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100000001100)
) lut_44_38 (
    .O(x44_y38),
    .I0(x42_y38),
    .I1(x42_y41),
    .I2(x41_y38),
    .I3(x42_y33)
);

(* keep, dont_touch *)
(* LOC = "X45/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111100010001)
) lut_45_38 (
    .O(x45_y38),
    .I0(x43_y36),
    .I1(x42_y40),
    .I2(x42_y34),
    .I3(x42_y33)
);

(* keep, dont_touch *)
(* LOC = "X46/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111010100011)
) lut_46_38 (
    .O(x46_y38),
    .I0(x44_y43),
    .I1(x44_y38),
    .I2(1'b0),
    .I3(x43_y37)
);

(* keep, dont_touch *)
(* LOC = "X47/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010011001100110)
) lut_47_38 (
    .O(x47_y38),
    .I0(x44_y40),
    .I1(x44_y38),
    .I2(x45_y39),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X48/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000100011000)
) lut_48_38 (
    .O(x48_y38),
    .I0(x46_y42),
    .I1(x45_y41),
    .I2(x46_y38),
    .I3(x45_y42)
);

(* keep, dont_touch *)
(* LOC = "X49/Y38" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110010110001)
) lut_49_38 (
    .O(x49_y38),
    .I0(x47_y33),
    .I1(x47_y33),
    .I2(x47_y34),
    .I3(x46_y41)
);

(* keep, dont_touch *)
(* LOC = "X0/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010100000101)
) lut_0_39 (
    .O(x0_y39),
    .I0(in1),
    .I1(in3),
    .I2(in3),
    .I3(in5)
);

(* keep, dont_touch *)
(* LOC = "X1/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111010110000)
) lut_1_39 (
    .O(x1_y39),
    .I0(in5),
    .I1(1'b0),
    .I2(in6),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X2/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010011100010)
) lut_2_39 (
    .O(x2_y39),
    .I0(in5),
    .I1(in8),
    .I2(in4),
    .I3(in4)
);

(* keep, dont_touch *)
(* LOC = "X3/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011001111001)
) lut_3_39 (
    .O(x3_y39),
    .I0(in5),
    .I1(x1_y41),
    .I2(in0),
    .I3(in5)
);

(* keep, dont_touch *)
(* LOC = "X4/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011001111001)
) lut_4_39 (
    .O(x4_y39),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X5/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011010001010)
) lut_5_39 (
    .O(x5_y39),
    .I0(1'b0),
    .I1(x2_y43),
    .I2(1'b0),
    .I3(x3_y42)
);

(* keep, dont_touch *)
(* LOC = "X6/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111011011100)
) lut_6_39 (
    .O(x6_y39),
    .I0(1'b0),
    .I1(x3_y35),
    .I2(1'b0),
    .I3(x4_y36)
);

(* keep, dont_touch *)
(* LOC = "X7/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100011110000)
) lut_7_39 (
    .O(x7_y39),
    .I0(x5_y39),
    .I1(x5_y44),
    .I2(x5_y41),
    .I3(x5_y38)
);

(* keep, dont_touch *)
(* LOC = "X8/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010010100011)
) lut_8_39 (
    .O(x8_y39),
    .I0(x6_y37),
    .I1(x6_y42),
    .I2(x6_y35),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X9/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010111110010)
) lut_9_39 (
    .O(x9_y39),
    .I0(x7_y37),
    .I1(x7_y44),
    .I2(x6_y35),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X10/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010011110111)
) lut_10_39 (
    .O(x10_y39),
    .I0(x7_y35),
    .I1(x8_y34),
    .I2(x7_y43),
    .I3(x8_y39)
);

(* keep, dont_touch *)
(* LOC = "X11/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011010100100)
) lut_11_39 (
    .O(x11_y39),
    .I0(1'b0),
    .I1(x8_y38),
    .I2(x8_y43),
    .I3(x8_y36)
);

(* keep, dont_touch *)
(* LOC = "X12/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101000101011)
) lut_12_39 (
    .O(x12_y39),
    .I0(x9_y38),
    .I1(x10_y44),
    .I2(1'b0),
    .I3(x10_y37)
);

(* keep, dont_touch *)
(* LOC = "X13/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110100011011)
) lut_13_39 (
    .O(x13_y39),
    .I0(1'b0),
    .I1(x11_y35),
    .I2(x10_y38),
    .I3(x11_y42)
);

(* keep, dont_touch *)
(* LOC = "X14/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000111010101)
) lut_14_39 (
    .O(x14_y39),
    .I0(x12_y37),
    .I1(1'b0),
    .I2(x12_y43),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X15/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000111110111)
) lut_15_39 (
    .O(x15_y39),
    .I0(x12_y36),
    .I1(x13_y38),
    .I2(x13_y37),
    .I3(x13_y42)
);

(* keep, dont_touch *)
(* LOC = "X16/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110111111111)
) lut_16_39 (
    .O(x16_y39),
    .I0(x13_y42),
    .I1(x14_y41),
    .I2(x14_y41),
    .I3(x14_y35)
);

(* keep, dont_touch *)
(* LOC = "X17/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010101110100)
) lut_17_39 (
    .O(x17_y39),
    .I0(1'b0),
    .I1(x15_y40),
    .I2(x14_y36),
    .I3(x14_y35)
);

(* keep, dont_touch *)
(* LOC = "X18/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000110111111)
) lut_18_39 (
    .O(x18_y39),
    .I0(x15_y40),
    .I1(1'b0),
    .I2(x15_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X19/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000110100100)
) lut_19_39 (
    .O(x19_y39),
    .I0(x17_y43),
    .I1(x16_y34),
    .I2(x16_y41),
    .I3(x16_y35)
);

(* keep, dont_touch *)
(* LOC = "X20/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101100111011)
) lut_20_39 (
    .O(x20_y39),
    .I0(x17_y38),
    .I1(x18_y34),
    .I2(x18_y38),
    .I3(x18_y44)
);

(* keep, dont_touch *)
(* LOC = "X21/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001101011001)
) lut_21_39 (
    .O(x21_y39),
    .I0(x19_y34),
    .I1(x18_y37),
    .I2(x18_y44),
    .I3(x18_y42)
);

(* keep, dont_touch *)
(* LOC = "X22/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001100111110)
) lut_22_39 (
    .O(x22_y39),
    .I0(1'b0),
    .I1(x20_y43),
    .I2(x19_y37),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X23/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101110100110)
) lut_23_39 (
    .O(x23_y39),
    .I0(x21_y41),
    .I1(x20_y44),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X24/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010010010110)
) lut_24_39 (
    .O(x24_y39),
    .I0(x22_y39),
    .I1(x21_y38),
    .I2(x22_y41),
    .I3(x21_y42)
);

(* keep, dont_touch *)
(* LOC = "X25/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100001001100)
) lut_25_39 (
    .O(x25_y39),
    .I0(x22_y39),
    .I1(x23_y35),
    .I2(x22_y38),
    .I3(x23_y39)
);

(* keep, dont_touch *)
(* LOC = "X26/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100111101111)
) lut_26_39 (
    .O(x26_y39),
    .I0(1'b0),
    .I1(x23_y38),
    .I2(x23_y36),
    .I3(x23_y37)
);

(* keep, dont_touch *)
(* LOC = "X27/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111101011101)
) lut_27_39 (
    .O(x27_y39),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x25_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X28/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100000110001)
) lut_28_39 (
    .O(x28_y39),
    .I0(x25_y42),
    .I1(x26_y36),
    .I2(1'b0),
    .I3(x25_y41)
);

(* keep, dont_touch *)
(* LOC = "X29/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101110000101)
) lut_29_39 (
    .O(x29_y39),
    .I0(1'b0),
    .I1(x27_y38),
    .I2(x27_y35),
    .I3(x27_y41)
);

(* keep, dont_touch *)
(* LOC = "X30/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010100100010)
) lut_30_39 (
    .O(x30_y39),
    .I0(x28_y38),
    .I1(x27_y35),
    .I2(x28_y40),
    .I3(x27_y35)
);

(* keep, dont_touch *)
(* LOC = "X31/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110101110000)
) lut_31_39 (
    .O(x31_y39),
    .I0(x29_y36),
    .I1(x29_y44),
    .I2(x29_y40),
    .I3(x28_y42)
);

(* keep, dont_touch *)
(* LOC = "X32/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101110100100)
) lut_32_39 (
    .O(x32_y39),
    .I0(x29_y42),
    .I1(x29_y36),
    .I2(1'b0),
    .I3(x30_y35)
);

(* keep, dont_touch *)
(* LOC = "X33/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101101001001)
) lut_33_39 (
    .O(x33_y39),
    .I0(x31_y39),
    .I1(x31_y41),
    .I2(x31_y42),
    .I3(x30_y38)
);

(* keep, dont_touch *)
(* LOC = "X34/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001111111111)
) lut_34_39 (
    .O(x34_y39),
    .I0(x32_y42),
    .I1(x31_y44),
    .I2(x31_y44),
    .I3(x31_y34)
);

(* keep, dont_touch *)
(* LOC = "X35/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000011000010)
) lut_35_39 (
    .O(x35_y39),
    .I0(x32_y43),
    .I1(x33_y34),
    .I2(x32_y42),
    .I3(x33_y41)
);

(* keep, dont_touch *)
(* LOC = "X36/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000110001100)
) lut_36_39 (
    .O(x36_y39),
    .I0(1'b0),
    .I1(x33_y37),
    .I2(x34_y40),
    .I3(x33_y42)
);

(* keep, dont_touch *)
(* LOC = "X37/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000110100110)
) lut_37_39 (
    .O(x37_y39),
    .I0(x34_y37),
    .I1(1'b0),
    .I2(x34_y38),
    .I3(x35_y41)
);

(* keep, dont_touch *)
(* LOC = "X38/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101111011110)
) lut_38_39 (
    .O(x38_y39),
    .I0(x35_y40),
    .I1(x35_y41),
    .I2(x36_y40),
    .I3(x35_y40)
);

(* keep, dont_touch *)
(* LOC = "X39/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011110111011)
) lut_39_39 (
    .O(x39_y39),
    .I0(x36_y37),
    .I1(x37_y41),
    .I2(x36_y43),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X40/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110110110100)
) lut_40_39 (
    .O(x40_y39),
    .I0(x37_y40),
    .I1(x38_y44),
    .I2(x38_y40),
    .I3(x37_y41)
);

(* keep, dont_touch *)
(* LOC = "X41/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000110111011)
) lut_41_39 (
    .O(x41_y39),
    .I0(x38_y40),
    .I1(x39_y37),
    .I2(x39_y35),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X42/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101010101010)
) lut_42_39 (
    .O(x42_y39),
    .I0(x39_y43),
    .I1(1'b0),
    .I2(x40_y39),
    .I3(x39_y39)
);

(* keep, dont_touch *)
(* LOC = "X43/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000001110010)
) lut_43_39 (
    .O(x43_y39),
    .I0(x41_y37),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x40_y37)
);

(* keep, dont_touch *)
(* LOC = "X44/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111111111001)
) lut_44_39 (
    .O(x44_y39),
    .I0(x42_y37),
    .I1(1'b0),
    .I2(x42_y34),
    .I3(x41_y36)
);

(* keep, dont_touch *)
(* LOC = "X45/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000101010011)
) lut_45_39 (
    .O(x45_y39),
    .I0(x43_y36),
    .I1(x42_y35),
    .I2(x42_y39),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X46/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000100100000)
) lut_46_39 (
    .O(x46_y39),
    .I0(1'b0),
    .I1(x43_y42),
    .I2(x44_y36),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X47/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101111110010)
) lut_47_39 (
    .O(x47_y39),
    .I0(x45_y35),
    .I1(x44_y43),
    .I2(1'b0),
    .I3(x45_y37)
);

(* keep, dont_touch *)
(* LOC = "X48/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000000001110)
) lut_48_39 (
    .O(x48_y39),
    .I0(x46_y39),
    .I1(x45_y36),
    .I2(x46_y39),
    .I3(x46_y37)
);

(* keep, dont_touch *)
(* LOC = "X49/Y39" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010111101101)
) lut_49_39 (
    .O(x49_y39),
    .I0(x47_y41),
    .I1(x47_y34),
    .I2(x47_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X0/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101010011100)
) lut_0_40 (
    .O(x0_y40),
    .I0(in8),
    .I1(in7),
    .I2(in1),
    .I3(in5)
);

(* keep, dont_touch *)
(* LOC = "X1/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100101111111)
) lut_1_40 (
    .O(x1_y40),
    .I0(in5),
    .I1(in1),
    .I2(in5),
    .I3(in7)
);

(* keep, dont_touch *)
(* LOC = "X2/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001001001010)
) lut_2_40 (
    .O(x2_y40),
    .I0(in5),
    .I1(in4),
    .I2(in6),
    .I3(in5)
);

(* keep, dont_touch *)
(* LOC = "X3/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111110101000)
) lut_3_40 (
    .O(x3_y40),
    .I0(1'b0),
    .I1(1'b0),
    .I2(in7),
    .I3(in2)
);

(* keep, dont_touch *)
(* LOC = "X4/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011100000001)
) lut_4_40 (
    .O(x4_y40),
    .I0(x2_y39),
    .I1(x1_y40),
    .I2(x2_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X5/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000101111101)
) lut_5_40 (
    .O(x5_y40),
    .I0(1'b0),
    .I1(x3_y39),
    .I2(1'b0),
    .I3(x2_y41)
);

(* keep, dont_touch *)
(* LOC = "X6/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010011101101)
) lut_6_40 (
    .O(x6_y40),
    .I0(x4_y41),
    .I1(x3_y37),
    .I2(x4_y38),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X7/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111010000010)
) lut_7_40 (
    .O(x7_y40),
    .I0(x4_y40),
    .I1(x4_y38),
    .I2(x5_y35),
    .I3(x4_y36)
);

(* keep, dont_touch *)
(* LOC = "X8/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101011101011)
) lut_8_40 (
    .O(x8_y40),
    .I0(x6_y43),
    .I1(x6_y44),
    .I2(x6_y38),
    .I3(x6_y40)
);

(* keep, dont_touch *)
(* LOC = "X9/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100101011001)
) lut_9_40 (
    .O(x9_y40),
    .I0(x7_y37),
    .I1(x6_y42),
    .I2(x6_y38),
    .I3(x6_y40)
);

(* keep, dont_touch *)
(* LOC = "X10/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001100011101)
) lut_10_40 (
    .O(x10_y40),
    .I0(x8_y42),
    .I1(1'b0),
    .I2(x8_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X11/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001011001011)
) lut_11_40 (
    .O(x11_y40),
    .I0(x8_y42),
    .I1(x8_y41),
    .I2(x8_y36),
    .I3(x9_y41)
);

(* keep, dont_touch *)
(* LOC = "X12/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001111000011)
) lut_12_40 (
    .O(x12_y40),
    .I0(x9_y37),
    .I1(1'b0),
    .I2(x10_y39),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X13/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110010110011)
) lut_13_40 (
    .O(x13_y40),
    .I0(x11_y44),
    .I1(x11_y40),
    .I2(x10_y36),
    .I3(x11_y42)
);

(* keep, dont_touch *)
(* LOC = "X14/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111010110011)
) lut_14_40 (
    .O(x14_y40),
    .I0(x12_y35),
    .I1(x11_y38),
    .I2(x12_y37),
    .I3(x12_y44)
);

(* keep, dont_touch *)
(* LOC = "X15/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111100111000)
) lut_15_40 (
    .O(x15_y40),
    .I0(1'b0),
    .I1(x12_y38),
    .I2(x13_y37),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X16/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101011001110)
) lut_16_40 (
    .O(x16_y40),
    .I0(x14_y39),
    .I1(x14_y45),
    .I2(x14_y37),
    .I3(x14_y42)
);

(* keep, dont_touch *)
(* LOC = "X17/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110111000111)
) lut_17_40 (
    .O(x17_y40),
    .I0(x14_y44),
    .I1(x14_y35),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X18/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010111001110)
) lut_18_40 (
    .O(x18_y40),
    .I0(x15_y41),
    .I1(x15_y43),
    .I2(x16_y38),
    .I3(x15_y36)
);

(* keep, dont_touch *)
(* LOC = "X19/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101101111111)
) lut_19_40 (
    .O(x19_y40),
    .I0(x16_y38),
    .I1(x16_y39),
    .I2(x16_y44),
    .I3(x16_y36)
);

(* keep, dont_touch *)
(* LOC = "X20/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100110110101)
) lut_20_40 (
    .O(x20_y40),
    .I0(x18_y43),
    .I1(x17_y37),
    .I2(x17_y43),
    .I3(x18_y39)
);

(* keep, dont_touch *)
(* LOC = "X21/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001000000100)
) lut_21_40 (
    .O(x21_y40),
    .I0(x18_y43),
    .I1(x19_y35),
    .I2(x19_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X22/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110010100100)
) lut_22_40 (
    .O(x22_y40),
    .I0(x19_y35),
    .I1(x20_y40),
    .I2(x20_y40),
    .I3(x19_y44)
);

(* keep, dont_touch *)
(* LOC = "X23/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101011100110)
) lut_23_40 (
    .O(x23_y40),
    .I0(x20_y44),
    .I1(x21_y39),
    .I2(x20_y41),
    .I3(x21_y41)
);

(* keep, dont_touch *)
(* LOC = "X24/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101110001000)
) lut_24_40 (
    .O(x24_y40),
    .I0(1'b0),
    .I1(x21_y40),
    .I2(x21_y43),
    .I3(x22_y45)
);

(* keep, dont_touch *)
(* LOC = "X25/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101101010100)
) lut_25_40 (
    .O(x25_y40),
    .I0(x22_y35),
    .I1(x22_y40),
    .I2(x23_y41),
    .I3(x22_y39)
);

(* keep, dont_touch *)
(* LOC = "X26/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001011110110)
) lut_26_40 (
    .O(x26_y40),
    .I0(1'b0),
    .I1(x24_y41),
    .I2(x24_y45),
    .I3(x24_y44)
);

(* keep, dont_touch *)
(* LOC = "X27/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111000011001)
) lut_27_40 (
    .O(x27_y40),
    .I0(x25_y35),
    .I1(x24_y38),
    .I2(1'b0),
    .I3(x24_y35)
);

(* keep, dont_touch *)
(* LOC = "X28/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101011011100)
) lut_28_40 (
    .O(x28_y40),
    .I0(x25_y45),
    .I1(x25_y35),
    .I2(x26_y42),
    .I3(x25_y36)
);

(* keep, dont_touch *)
(* LOC = "X29/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000011000101)
) lut_29_40 (
    .O(x29_y40),
    .I0(x27_y36),
    .I1(x26_y36),
    .I2(x26_y40),
    .I3(x27_y38)
);

(* keep, dont_touch *)
(* LOC = "X30/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110000111000)
) lut_30_40 (
    .O(x30_y40),
    .I0(x28_y41),
    .I1(x27_y36),
    .I2(x27_y35),
    .I3(x27_y36)
);

(* keep, dont_touch *)
(* LOC = "X31/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110010110000)
) lut_31_40 (
    .O(x31_y40),
    .I0(x28_y37),
    .I1(x28_y38),
    .I2(x29_y44),
    .I3(x29_y37)
);

(* keep, dont_touch *)
(* LOC = "X32/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010101001111)
) lut_32_40 (
    .O(x32_y40),
    .I0(x29_y37),
    .I1(x29_y38),
    .I2(x29_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X33/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011110110011)
) lut_33_40 (
    .O(x33_y40),
    .I0(x31_y35),
    .I1(x30_y44),
    .I2(x31_y36),
    .I3(x31_y42)
);

(* keep, dont_touch *)
(* LOC = "X34/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001101111101)
) lut_34_40 (
    .O(x34_y40),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x32_y37),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X35/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001101101001)
) lut_35_40 (
    .O(x35_y40),
    .I0(x33_y40),
    .I1(1'b0),
    .I2(x33_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X36/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100101001011)
) lut_36_40 (
    .O(x36_y40),
    .I0(x33_y36),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x34_y43)
);

(* keep, dont_touch *)
(* LOC = "X37/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001001100001)
) lut_37_40 (
    .O(x37_y40),
    .I0(x35_y35),
    .I1(1'b0),
    .I2(x34_y43),
    .I3(x35_y35)
);

(* keep, dont_touch *)
(* LOC = "X38/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011010111111)
) lut_38_40 (
    .O(x38_y40),
    .I0(x36_y43),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X39/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110100001000)
) lut_39_40 (
    .O(x39_y40),
    .I0(1'b0),
    .I1(x37_y39),
    .I2(x36_y44),
    .I3(x37_y36)
);

(* keep, dont_touch *)
(* LOC = "X40/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111011010101)
) lut_40_40 (
    .O(x40_y40),
    .I0(x37_y42),
    .I1(1'b0),
    .I2(x37_y41),
    .I3(x37_y38)
);

(* keep, dont_touch *)
(* LOC = "X41/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011011011011)
) lut_41_40 (
    .O(x41_y40),
    .I0(x39_y36),
    .I1(1'b0),
    .I2(x38_y35),
    .I3(x38_y36)
);

(* keep, dont_touch *)
(* LOC = "X42/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111011010101)
) lut_42_40 (
    .O(x42_y40),
    .I0(x40_y37),
    .I1(x39_y43),
    .I2(x40_y40),
    .I3(x40_y36)
);

(* keep, dont_touch *)
(* LOC = "X43/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110000111010)
) lut_43_40 (
    .O(x43_y40),
    .I0(x41_y36),
    .I1(x40_y38),
    .I2(x40_y41),
    .I3(x40_y35)
);

(* keep, dont_touch *)
(* LOC = "X44/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101001111100)
) lut_44_40 (
    .O(x44_y40),
    .I0(x41_y42),
    .I1(1'b0),
    .I2(x41_y45),
    .I3(x42_y41)
);

(* keep, dont_touch *)
(* LOC = "X45/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110010100111)
) lut_45_40 (
    .O(x45_y40),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x42_y45),
    .I3(x43_y41)
);

(* keep, dont_touch *)
(* LOC = "X46/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001111101111)
) lut_46_40 (
    .O(x46_y40),
    .I0(x44_y39),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x44_y36)
);

(* keep, dont_touch *)
(* LOC = "X47/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000100000101)
) lut_47_40 (
    .O(x47_y40),
    .I0(x44_y39),
    .I1(x45_y42),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X48/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101010111100)
) lut_48_40 (
    .O(x48_y40),
    .I0(1'b0),
    .I1(x45_y40),
    .I2(x45_y35),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X49/Y40" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100101101000)
) lut_49_40 (
    .O(x49_y40),
    .I0(1'b0),
    .I1(x47_y35),
    .I2(x46_y36),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X0/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100101011110)
) lut_0_41 (
    .O(x0_y41),
    .I0(in7),
    .I1(in8),
    .I2(in7),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X1/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000010001000)
) lut_1_41 (
    .O(x1_y41),
    .I0(1'b0),
    .I1(1'b0),
    .I2(in1),
    .I3(in2)
);

(* keep, dont_touch *)
(* LOC = "X2/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101111010000)
) lut_2_41 (
    .O(x2_y41),
    .I0(1'b0),
    .I1(in2),
    .I2(in0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X3/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101011101010)
) lut_3_41 (
    .O(x3_y41),
    .I0(x1_y42),
    .I1(in0),
    .I2(in6),
    .I3(in6)
);

(* keep, dont_touch *)
(* LOC = "X4/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111001010110)
) lut_4_41 (
    .O(x4_y41),
    .I0(x1_y37),
    .I1(x1_y42),
    .I2(x2_y41),
    .I3(x1_y40)
);

(* keep, dont_touch *)
(* LOC = "X5/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011011110010)
) lut_5_41 (
    .O(x5_y41),
    .I0(x2_y46),
    .I1(x2_y36),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X6/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010111110101)
) lut_6_41 (
    .O(x6_y41),
    .I0(x4_y44),
    .I1(1'b0),
    .I2(x4_y41),
    .I3(x3_y36)
);

(* keep, dont_touch *)
(* LOC = "X7/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101110111101010)
) lut_7_41 (
    .O(x7_y41),
    .I0(x4_y46),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x5_y46)
);

(* keep, dont_touch *)
(* LOC = "X8/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000101110010)
) lut_8_41 (
    .O(x8_y41),
    .I0(x6_y43),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X9/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011111010111)
) lut_9_41 (
    .O(x9_y41),
    .I0(x6_y41),
    .I1(x6_y46),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X10/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010001000010)
) lut_10_41 (
    .O(x10_y41),
    .I0(x7_y41),
    .I1(x8_y42),
    .I2(1'b0),
    .I3(x8_y40)
);

(* keep, dont_touch *)
(* LOC = "X11/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010001010010)
) lut_11_41 (
    .O(x11_y41),
    .I0(x9_y40),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x9_y40)
);

(* keep, dont_touch *)
(* LOC = "X12/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010101110100)
) lut_12_41 (
    .O(x12_y41),
    .I0(1'b0),
    .I1(x10_y46),
    .I2(x9_y42),
    .I3(x9_y42)
);

(* keep, dont_touch *)
(* LOC = "X13/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110000000101)
) lut_13_41 (
    .O(x13_y41),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x10_y44),
    .I3(x10_y41)
);

(* keep, dont_touch *)
(* LOC = "X14/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011010110110)
) lut_14_41 (
    .O(x14_y41),
    .I0(x12_y43),
    .I1(x11_y40),
    .I2(x11_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X15/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010010011000)
) lut_15_41 (
    .O(x15_y41),
    .I0(x13_y39),
    .I1(x13_y44),
    .I2(1'b0),
    .I3(x12_y37)
);

(* keep, dont_touch *)
(* LOC = "X16/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000100100101)
) lut_16_41 (
    .O(x16_y41),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x14_y39),
    .I3(x14_y45)
);

(* keep, dont_touch *)
(* LOC = "X17/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011011111011)
) lut_17_41 (
    .O(x17_y41),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x15_y40)
);

(* keep, dont_touch *)
(* LOC = "X18/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000101100101)
) lut_18_41 (
    .O(x18_y41),
    .I0(x15_y38),
    .I1(1'b0),
    .I2(x16_y38),
    .I3(x16_y41)
);

(* keep, dont_touch *)
(* LOC = "X19/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011001001001)
) lut_19_41 (
    .O(x19_y41),
    .I0(x16_y41),
    .I1(x17_y41),
    .I2(x16_y41),
    .I3(x16_y36)
);

(* keep, dont_touch *)
(* LOC = "X20/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001000010101)
) lut_20_41 (
    .O(x20_y41),
    .I0(x18_y44),
    .I1(x18_y43),
    .I2(x18_y45),
    .I3(x18_y36)
);

(* keep, dont_touch *)
(* LOC = "X21/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011001111110)
) lut_21_41 (
    .O(x21_y41),
    .I0(x19_y46),
    .I1(x19_y45),
    .I2(x19_y40),
    .I3(x18_y40)
);

(* keep, dont_touch *)
(* LOC = "X22/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101101001111)
) lut_22_41 (
    .O(x22_y41),
    .I0(x20_y45),
    .I1(x19_y40),
    .I2(x20_y43),
    .I3(x19_y44)
);

(* keep, dont_touch *)
(* LOC = "X23/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000010001001)
) lut_23_41 (
    .O(x23_y41),
    .I0(x20_y46),
    .I1(x21_y41),
    .I2(x21_y41),
    .I3(x21_y44)
);

(* keep, dont_touch *)
(* LOC = "X24/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110100000110)
) lut_24_41 (
    .O(x24_y41),
    .I0(1'b0),
    .I1(x21_y46),
    .I2(1'b0),
    .I3(x21_y45)
);

(* keep, dont_touch *)
(* LOC = "X25/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010011000010)
) lut_25_41 (
    .O(x25_y41),
    .I0(x22_y37),
    .I1(x23_y37),
    .I2(x22_y43),
    .I3(x22_y37)
);

(* keep, dont_touch *)
(* LOC = "X26/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100101100111)
) lut_26_41 (
    .O(x26_y41),
    .I0(x24_y38),
    .I1(x24_y42),
    .I2(x24_y42),
    .I3(x23_y41)
);

(* keep, dont_touch *)
(* LOC = "X27/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011000001110)
) lut_27_41 (
    .O(x27_y41),
    .I0(1'b0),
    .I1(x25_y46),
    .I2(x25_y42),
    .I3(x24_y36)
);

(* keep, dont_touch *)
(* LOC = "X28/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001000101111)
) lut_28_41 (
    .O(x28_y41),
    .I0(x25_y41),
    .I1(x26_y41),
    .I2(1'b0),
    .I3(x26_y41)
);

(* keep, dont_touch *)
(* LOC = "X29/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111000011110)
) lut_29_41 (
    .O(x29_y41),
    .I0(x27_y45),
    .I1(1'b0),
    .I2(x27_y41),
    .I3(x26_y44)
);

(* keep, dont_touch *)
(* LOC = "X30/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011010111110)
) lut_30_41 (
    .O(x30_y41),
    .I0(1'b0),
    .I1(x27_y44),
    .I2(x27_y43),
    .I3(x28_y46)
);

(* keep, dont_touch *)
(* LOC = "X31/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111000101001)
) lut_31_41 (
    .O(x31_y41),
    .I0(1'b0),
    .I1(x29_y38),
    .I2(x29_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X32/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101101011100)
) lut_32_41 (
    .O(x32_y41),
    .I0(x29_y40),
    .I1(x30_y36),
    .I2(x30_y45),
    .I3(x29_y46)
);

(* keep, dont_touch *)
(* LOC = "X33/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101001001101)
) lut_33_41 (
    .O(x33_y41),
    .I0(x30_y39),
    .I1(x31_y46),
    .I2(1'b0),
    .I3(x31_y46)
);

(* keep, dont_touch *)
(* LOC = "X34/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011010110111)
) lut_34_41 (
    .O(x34_y41),
    .I0(1'b0),
    .I1(x31_y45),
    .I2(x31_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X35/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000100011000)
) lut_35_41 (
    .O(x35_y41),
    .I0(x33_y38),
    .I1(x32_y41),
    .I2(x32_y45),
    .I3(x32_y45)
);

(* keep, dont_touch *)
(* LOC = "X36/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111001010111)
) lut_36_41 (
    .O(x36_y41),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x33_y46),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X37/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100011010011)
) lut_37_41 (
    .O(x37_y41),
    .I0(x34_y42),
    .I1(1'b0),
    .I2(x35_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X38/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000000111100)
) lut_38_41 (
    .O(x38_y41),
    .I0(1'b0),
    .I1(x36_y36),
    .I2(1'b0),
    .I3(x35_y46)
);

(* keep, dont_touch *)
(* LOC = "X39/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101000111010)
) lut_39_41 (
    .O(x39_y41),
    .I0(x37_y45),
    .I1(x36_y38),
    .I2(x37_y44),
    .I3(x36_y42)
);

(* keep, dont_touch *)
(* LOC = "X40/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010010110001)
) lut_40_41 (
    .O(x40_y41),
    .I0(x38_y36),
    .I1(x37_y41),
    .I2(x37_y46),
    .I3(x38_y36)
);

(* keep, dont_touch *)
(* LOC = "X41/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011110111001)
) lut_41_41 (
    .O(x41_y41),
    .I0(1'b0),
    .I1(x39_y41),
    .I2(x38_y39),
    .I3(x39_y38)
);

(* keep, dont_touch *)
(* LOC = "X42/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111000100001)
) lut_42_41 (
    .O(x42_y41),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x39_y42),
    .I3(x40_y42)
);

(* keep, dont_touch *)
(* LOC = "X43/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010110000110)
) lut_43_41 (
    .O(x43_y41),
    .I0(1'b0),
    .I1(x41_y44),
    .I2(x41_y36),
    .I3(x40_y40)
);

(* keep, dont_touch *)
(* LOC = "X44/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000010100001)
) lut_44_41 (
    .O(x44_y41),
    .I0(1'b0),
    .I1(x41_y44),
    .I2(x42_y38),
    .I3(x42_y37)
);

(* keep, dont_touch *)
(* LOC = "X45/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011001110001)
) lut_45_41 (
    .O(x45_y41),
    .I0(x43_y46),
    .I1(x42_y36),
    .I2(1'b0),
    .I3(x42_y40)
);

(* keep, dont_touch *)
(* LOC = "X46/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001000110011)
) lut_46_41 (
    .O(x46_y41),
    .I0(x44_y41),
    .I1(x44_y46),
    .I2(1'b0),
    .I3(x44_y42)
);

(* keep, dont_touch *)
(* LOC = "X47/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110101010100)
) lut_47_41 (
    .O(x47_y41),
    .I0(x45_y41),
    .I1(x44_y39),
    .I2(x44_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X48/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111110110101100)
) lut_48_41 (
    .O(x48_y41),
    .I0(x45_y38),
    .I1(1'b0),
    .I2(x46_y44),
    .I3(x46_y38)
);

(* keep, dont_touch *)
(* LOC = "X49/Y41" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001101100100)
) lut_49_41 (
    .O(x49_y41),
    .I0(x47_y39),
    .I1(x47_y41),
    .I2(x47_y37),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X0/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110100101110)
) lut_0_42 (
    .O(x0_y42),
    .I0(in3),
    .I1(1'b0),
    .I2(in6),
    .I3(in8)
);

(* keep, dont_touch *)
(* LOC = "X1/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101111101101)
) lut_1_42 (
    .O(x1_y42),
    .I0(in1),
    .I1(in3),
    .I2(in3),
    .I3(in9)
);

(* keep, dont_touch *)
(* LOC = "X2/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111011110010)
) lut_2_42 (
    .O(x2_y42),
    .I0(in7),
    .I1(in3),
    .I2(in3),
    .I3(in3)
);

(* keep, dont_touch *)
(* LOC = "X3/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010010001101)
) lut_3_42 (
    .O(x3_y42),
    .I0(in4),
    .I1(x1_y44),
    .I2(in0),
    .I3(x1_y40)
);

(* keep, dont_touch *)
(* LOC = "X4/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111101000000)
) lut_4_42 (
    .O(x4_y42),
    .I0(x1_y38),
    .I1(1'b0),
    .I2(x1_y47),
    .I3(x2_y47)
);

(* keep, dont_touch *)
(* LOC = "X5/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110001110101)
) lut_5_42 (
    .O(x5_y42),
    .I0(x3_y45),
    .I1(x2_y37),
    .I2(1'b0),
    .I3(x2_y43)
);

(* keep, dont_touch *)
(* LOC = "X6/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101111011010)
) lut_6_42 (
    .O(x6_y42),
    .I0(x4_y37),
    .I1(x4_y41),
    .I2(x3_y43),
    .I3(x4_y38)
);

(* keep, dont_touch *)
(* LOC = "X7/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000100010101)
) lut_7_42 (
    .O(x7_y42),
    .I0(x4_y47),
    .I1(1'b0),
    .I2(x4_y46),
    .I3(x5_y39)
);

(* keep, dont_touch *)
(* LOC = "X8/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011010110001)
) lut_8_42 (
    .O(x8_y42),
    .I0(x6_y46),
    .I1(x6_y40),
    .I2(x5_y40),
    .I3(x5_y40)
);

(* keep, dont_touch *)
(* LOC = "X9/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011001001000)
) lut_9_42 (
    .O(x9_y42),
    .I0(x7_y38),
    .I1(1'b0),
    .I2(x5_y40),
    .I3(x5_y40)
);

(* keep, dont_touch *)
(* LOC = "X10/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011111001000)
) lut_10_42 (
    .O(x10_y42),
    .I0(x8_y45),
    .I1(x7_y37),
    .I2(x7_y41),
    .I3(x8_y40)
);

(* keep, dont_touch *)
(* LOC = "X11/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110001011110111)
) lut_11_42 (
    .O(x11_y42),
    .I0(x9_y45),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x8_y39)
);

(* keep, dont_touch *)
(* LOC = "X12/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000011011111)
) lut_12_42 (
    .O(x12_y42),
    .I0(1'b0),
    .I1(x9_y42),
    .I2(x10_y37),
    .I3(x10_y44)
);

(* keep, dont_touch *)
(* LOC = "X13/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110011111001)
) lut_13_42 (
    .O(x13_y42),
    .I0(x10_y41),
    .I1(x10_y45),
    .I2(x11_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X14/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011111100100)
) lut_14_42 (
    .O(x14_y42),
    .I0(x11_y45),
    .I1(x12_y42),
    .I2(1'b0),
    .I3(x12_y37)
);

(* keep, dont_touch *)
(* LOC = "X15/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110111110000)
) lut_15_42 (
    .O(x15_y42),
    .I0(x12_y38),
    .I1(x13_y42),
    .I2(x12_y40),
    .I3(x12_y39)
);

(* keep, dont_touch *)
(* LOC = "X16/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110010100110)
) lut_16_42 (
    .O(x16_y42),
    .I0(1'b0),
    .I1(x14_y39),
    .I2(x13_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X17/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011000111100)
) lut_17_42 (
    .O(x17_y42),
    .I0(x14_y45),
    .I1(1'b0),
    .I2(x15_y39),
    .I3(x15_y38)
);

(* keep, dont_touch *)
(* LOC = "X18/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011100101111)
) lut_18_42 (
    .O(x18_y42),
    .I0(x15_y41),
    .I1(x15_y39),
    .I2(x15_y37),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X19/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000111011101)
) lut_19_42 (
    .O(x19_y42),
    .I0(x16_y47),
    .I1(1'b0),
    .I2(x17_y42),
    .I3(x17_y38)
);

(* keep, dont_touch *)
(* LOC = "X20/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010110011100)
) lut_20_42 (
    .O(x20_y42),
    .I0(x17_y39),
    .I1(x17_y38),
    .I2(x17_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X21/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110110000101)
) lut_21_42 (
    .O(x21_y42),
    .I0(1'b0),
    .I1(x18_y43),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X22/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101010000001101)
) lut_22_42 (
    .O(x22_y42),
    .I0(1'b0),
    .I1(x19_y38),
    .I2(1'b0),
    .I3(x19_y45)
);

(* keep, dont_touch *)
(* LOC = "X23/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001101001110)
) lut_23_42 (
    .O(x23_y42),
    .I0(x21_y43),
    .I1(x21_y37),
    .I2(x20_y37),
    .I3(x20_y47)
);

(* keep, dont_touch *)
(* LOC = "X24/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101100111100)
) lut_24_42 (
    .O(x24_y42),
    .I0(x22_y43),
    .I1(x21_y47),
    .I2(x22_y39),
    .I3(x21_y37)
);

(* keep, dont_touch *)
(* LOC = "X25/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010101011010)
) lut_25_42 (
    .O(x25_y42),
    .I0(1'b0),
    .I1(x22_y45),
    .I2(x23_y42),
    .I3(x23_y47)
);

(* keep, dont_touch *)
(* LOC = "X26/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100100100010)
) lut_26_42 (
    .O(x26_y42),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x24_y38),
    .I3(x24_y37)
);

(* keep, dont_touch *)
(* LOC = "X27/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011001110001)
) lut_27_42 (
    .O(x27_y42),
    .I0(1'b0),
    .I1(x24_y47),
    .I2(x24_y43),
    .I3(x24_y39)
);

(* keep, dont_touch *)
(* LOC = "X28/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111010010111)
) lut_28_42 (
    .O(x28_y42),
    .I0(1'b0),
    .I1(x26_y40),
    .I2(x25_y46),
    .I3(x25_y46)
);

(* keep, dont_touch *)
(* LOC = "X29/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000011110111)
) lut_29_42 (
    .O(x29_y42),
    .I0(1'b0),
    .I1(x27_y45),
    .I2(x26_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X30/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101100100110)
) lut_30_42 (
    .O(x30_y42),
    .I0(x28_y46),
    .I1(x27_y40),
    .I2(x27_y38),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X31/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101011101011)
) lut_31_42 (
    .O(x31_y42),
    .I0(x28_y47),
    .I1(x29_y40),
    .I2(x29_y40),
    .I3(x29_y40)
);

(* keep, dont_touch *)
(* LOC = "X32/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110110110010)
) lut_32_42 (
    .O(x32_y42),
    .I0(x30_y38),
    .I1(x29_y38),
    .I2(x29_y38),
    .I3(x29_y41)
);

(* keep, dont_touch *)
(* LOC = "X33/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101010100111)
) lut_33_42 (
    .O(x33_y42),
    .I0(x31_y39),
    .I1(x31_y39),
    .I2(x30_y44),
    .I3(x31_y46)
);

(* keep, dont_touch *)
(* LOC = "X34/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101010010110)
) lut_34_42 (
    .O(x34_y42),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X35/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110111010010)
) lut_35_42 (
    .O(x35_y42),
    .I0(x32_y44),
    .I1(x33_y46),
    .I2(x32_y40),
    .I3(x33_y37)
);

(* keep, dont_touch *)
(* LOC = "X36/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000100111001)
) lut_36_42 (
    .O(x36_y42),
    .I0(1'b0),
    .I1(x34_y47),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X37/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000011100000)
) lut_37_42 (
    .O(x37_y42),
    .I0(x35_y41),
    .I1(x34_y41),
    .I2(x35_y37),
    .I3(x35_y39)
);

(* keep, dont_touch *)
(* LOC = "X38/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101101000100)
) lut_38_42 (
    .O(x38_y42),
    .I0(x36_y44),
    .I1(x35_y39),
    .I2(x36_y41),
    .I3(x36_y42)
);

(* keep, dont_touch *)
(* LOC = "X39/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110011101001)
) lut_39_42 (
    .O(x39_y42),
    .I0(x36_y40),
    .I1(x37_y45),
    .I2(x37_y37),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X40/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001110010100101)
) lut_40_42 (
    .O(x40_y42),
    .I0(x38_y47),
    .I1(1'b0),
    .I2(x37_y46),
    .I3(x37_y38)
);

(* keep, dont_touch *)
(* LOC = "X41/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010011010100)
) lut_41_42 (
    .O(x41_y42),
    .I0(x38_y44),
    .I1(x38_y37),
    .I2(x39_y38),
    .I3(x39_y44)
);

(* keep, dont_touch *)
(* LOC = "X42/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111100111011)
) lut_42_42 (
    .O(x42_y42),
    .I0(x40_y40),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x40_y40)
);

(* keep, dont_touch *)
(* LOC = "X43/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010101110101)
) lut_43_42 (
    .O(x43_y42),
    .I0(x41_y40),
    .I1(x41_y45),
    .I2(1'b0),
    .I3(x40_y40)
);

(* keep, dont_touch *)
(* LOC = "X44/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001111111100)
) lut_44_42 (
    .O(x44_y42),
    .I0(1'b0),
    .I1(x42_y41),
    .I2(1'b0),
    .I3(x42_y44)
);

(* keep, dont_touch *)
(* LOC = "X45/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011011000111)
) lut_45_42 (
    .O(x45_y42),
    .I0(x42_y46),
    .I1(x42_y37),
    .I2(x43_y38),
    .I3(x42_y38)
);

(* keep, dont_touch *)
(* LOC = "X46/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010000001100)
) lut_46_42 (
    .O(x46_y42),
    .I0(x44_y37),
    .I1(x44_y37),
    .I2(x44_y46),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X47/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001010101100)
) lut_47_42 (
    .O(x47_y42),
    .I0(x44_y45),
    .I1(x45_y45),
    .I2(x44_y46),
    .I3(x45_y40)
);

(* keep, dont_touch *)
(* LOC = "X48/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001101011001)
) lut_48_42 (
    .O(x48_y42),
    .I0(x45_y41),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X49/Y42" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101001011110)
) lut_49_42 (
    .O(x49_y42),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x46_y45),
    .I3(x46_y37)
);

(* keep, dont_touch *)
(* LOC = "X0/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011101101100)
) lut_0_43 (
    .O(x0_y43),
    .I0(in9),
    .I1(in8),
    .I2(in7),
    .I3(in0)
);

(* keep, dont_touch *)
(* LOC = "X1/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011010011010)
) lut_1_43 (
    .O(x1_y43),
    .I0(in0),
    .I1(in4),
    .I2(in7),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X2/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111110111111)
) lut_2_43 (
    .O(x2_y43),
    .I0(1'b0),
    .I1(in2),
    .I2(in1),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X3/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101111100110)
) lut_3_43 (
    .O(x3_y43),
    .I0(in2),
    .I1(in4),
    .I2(in6),
    .I3(x1_y44)
);

(* keep, dont_touch *)
(* LOC = "X4/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010001001000)
) lut_4_43 (
    .O(x4_y43),
    .I0(x1_y43),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x1_y46)
);

(* keep, dont_touch *)
(* LOC = "X5/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010111001111)
) lut_5_43 (
    .O(x5_y43),
    .I0(x3_y48),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x2_y42)
);

(* keep, dont_touch *)
(* LOC = "X6/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011101010101)
) lut_6_43 (
    .O(x6_y43),
    .I0(x3_y38),
    .I1(x3_y40),
    .I2(x4_y39),
    .I3(x4_y45)
);

(* keep, dont_touch *)
(* LOC = "X7/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111010100111)
) lut_7_43 (
    .O(x7_y43),
    .I0(x5_y41),
    .I1(x5_y38),
    .I2(x4_y43),
    .I3(x4_y43)
);

(* keep, dont_touch *)
(* LOC = "X8/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001111011101)
) lut_8_43 (
    .O(x8_y43),
    .I0(x5_y47),
    .I1(x5_y41),
    .I2(x5_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X9/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000100100010)
) lut_9_43 (
    .O(x9_y43),
    .I0(x7_y48),
    .I1(x6_y42),
    .I2(x5_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X10/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101111110011)
) lut_10_43 (
    .O(x10_y43),
    .I0(x7_y47),
    .I1(x7_y40),
    .I2(x7_y48),
    .I3(x8_y43)
);

(* keep, dont_touch *)
(* LOC = "X11/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100010101111)
) lut_11_43 (
    .O(x11_y43),
    .I0(1'b0),
    .I1(x9_y48),
    .I2(x8_y42),
    .I3(x8_y39)
);

(* keep, dont_touch *)
(* LOC = "X12/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010111000100010)
) lut_12_43 (
    .O(x12_y43),
    .I0(x10_y47),
    .I1(x9_y45),
    .I2(x10_y44),
    .I3(x10_y45)
);

(* keep, dont_touch *)
(* LOC = "X13/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111000101110)
) lut_13_43 (
    .O(x13_y43),
    .I0(1'b0),
    .I1(x11_y48),
    .I2(x10_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X14/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100001010101)
) lut_14_43 (
    .O(x14_y43),
    .I0(x12_y38),
    .I1(x11_y46),
    .I2(x11_y44),
    .I3(x12_y46)
);

(* keep, dont_touch *)
(* LOC = "X15/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101001001101)
) lut_15_43 (
    .O(x15_y43),
    .I0(1'b0),
    .I1(x13_y48),
    .I2(x13_y44),
    .I3(x13_y48)
);

(* keep, dont_touch *)
(* LOC = "X16/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001001111010)
) lut_16_43 (
    .O(x16_y43),
    .I0(x14_y42),
    .I1(x13_y44),
    .I2(x14_y44),
    .I3(x13_y39)
);

(* keep, dont_touch *)
(* LOC = "X17/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100101111000)
) lut_17_43 (
    .O(x17_y43),
    .I0(x15_y45),
    .I1(x14_y42),
    .I2(x14_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X18/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101101101000)
) lut_18_43 (
    .O(x18_y43),
    .I0(x16_y48),
    .I1(x15_y46),
    .I2(x16_y44),
    .I3(x16_y46)
);

(* keep, dont_touch *)
(* LOC = "X19/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110001101010101)
) lut_19_43 (
    .O(x19_y43),
    .I0(x17_y40),
    .I1(x17_y38),
    .I2(x16_y38),
    .I3(x17_y39)
);

(* keep, dont_touch *)
(* LOC = "X20/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101010110011)
) lut_20_43 (
    .O(x20_y43),
    .I0(x18_y46),
    .I1(x18_y38),
    .I2(x18_y39),
    .I3(x17_y46)
);

(* keep, dont_touch *)
(* LOC = "X21/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011000010111)
) lut_21_43 (
    .O(x21_y43),
    .I0(x19_y44),
    .I1(x19_y39),
    .I2(1'b0),
    .I3(x19_y43)
);

(* keep, dont_touch *)
(* LOC = "X22/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011111011101)
) lut_22_43 (
    .O(x22_y43),
    .I0(x19_y43),
    .I1(x20_y46),
    .I2(x20_y40),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X23/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111010010010)
) lut_23_43 (
    .O(x23_y43),
    .I0(1'b0),
    .I1(x21_y44),
    .I2(x20_y40),
    .I3(x21_y38)
);

(* keep, dont_touch *)
(* LOC = "X24/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110000110110)
) lut_24_43 (
    .O(x24_y43),
    .I0(x21_y47),
    .I1(x21_y47),
    .I2(x21_y43),
    .I3(x22_y47)
);

(* keep, dont_touch *)
(* LOC = "X25/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101110101100)
) lut_25_43 (
    .O(x25_y43),
    .I0(x23_y45),
    .I1(x23_y48),
    .I2(1'b0),
    .I3(x23_y43)
);

(* keep, dont_touch *)
(* LOC = "X26/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001111111101001)
) lut_26_43 (
    .O(x26_y43),
    .I0(x24_y45),
    .I1(1'b0),
    .I2(x24_y44),
    .I3(x24_y38)
);

(* keep, dont_touch *)
(* LOC = "X27/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101000001100)
) lut_27_43 (
    .O(x27_y43),
    .I0(x25_y43),
    .I1(x24_y43),
    .I2(x25_y39),
    .I3(x24_y44)
);

(* keep, dont_touch *)
(* LOC = "X28/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011011011111)
) lut_28_43 (
    .O(x28_y43),
    .I0(x25_y38),
    .I1(x26_y39),
    .I2(1'b0),
    .I3(x26_y38)
);

(* keep, dont_touch *)
(* LOC = "X29/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001111010110)
) lut_29_43 (
    .O(x29_y43),
    .I0(x27_y46),
    .I1(x27_y46),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X30/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001001001100)
) lut_30_43 (
    .O(x30_y43),
    .I0(x28_y47),
    .I1(x28_y38),
    .I2(x27_y42),
    .I3(x27_y42)
);

(* keep, dont_touch *)
(* LOC = "X31/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001000101001)
) lut_31_43 (
    .O(x31_y43),
    .I0(x28_y42),
    .I1(x28_y46),
    .I2(x29_y42),
    .I3(x28_y39)
);

(* keep, dont_touch *)
(* LOC = "X32/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100110101101)
) lut_32_43 (
    .O(x32_y43),
    .I0(1'b0),
    .I1(x30_y47),
    .I2(x29_y38),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X33/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100111101111)
) lut_33_43 (
    .O(x33_y43),
    .I0(x30_y48),
    .I1(1'b0),
    .I2(x30_y42),
    .I3(x30_y41)
);

(* keep, dont_touch *)
(* LOC = "X34/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101000001010)
) lut_34_43 (
    .O(x34_y43),
    .I0(x32_y39),
    .I1(1'b0),
    .I2(x31_y41),
    .I3(x32_y38)
);

(* keep, dont_touch *)
(* LOC = "X35/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100111100011101)
) lut_35_43 (
    .O(x35_y43),
    .I0(1'b0),
    .I1(x32_y46),
    .I2(x33_y45),
    .I3(x32_y42)
);

(* keep, dont_touch *)
(* LOC = "X36/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100101100010)
) lut_36_43 (
    .O(x36_y43),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x34_y43),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X37/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010100100000)
) lut_37_43 (
    .O(x37_y43),
    .I0(x35_y38),
    .I1(x35_y43),
    .I2(x34_y41),
    .I3(x35_y40)
);

(* keep, dont_touch *)
(* LOC = "X38/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010011000011)
) lut_38_43 (
    .O(x38_y43),
    .I0(x36_y42),
    .I1(1'b0),
    .I2(x36_y44),
    .I3(x35_y46)
);

(* keep, dont_touch *)
(* LOC = "X39/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011100010100)
) lut_39_43 (
    .O(x39_y43),
    .I0(x36_y40),
    .I1(x37_y43),
    .I2(x36_y39),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X40/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001110110110)
) lut_40_43 (
    .O(x40_y43),
    .I0(x37_y38),
    .I1(1'b0),
    .I2(x37_y40),
    .I3(x38_y47)
);

(* keep, dont_touch *)
(* LOC = "X41/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100100111011)
) lut_41_43 (
    .O(x41_y43),
    .I0(1'b0),
    .I1(x38_y40),
    .I2(1'b0),
    .I3(x38_y38)
);

(* keep, dont_touch *)
(* LOC = "X42/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001101001001)
) lut_42_43 (
    .O(x42_y43),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x39_y45),
    .I3(x40_y43)
);

(* keep, dont_touch *)
(* LOC = "X43/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111110111100)
) lut_43_43 (
    .O(x43_y43),
    .I0(x40_y42),
    .I1(x41_y38),
    .I2(x40_y39),
    .I3(x41_y47)
);

(* keep, dont_touch *)
(* LOC = "X44/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011110111110)
) lut_44_43 (
    .O(x44_y43),
    .I0(1'b0),
    .I1(x42_y38),
    .I2(x41_y47),
    .I3(x41_y46)
);

(* keep, dont_touch *)
(* LOC = "X45/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100110010101010)
) lut_45_43 (
    .O(x45_y43),
    .I0(x42_y45),
    .I1(x43_y39),
    .I2(x43_y41),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X46/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100011000100)
) lut_46_43 (
    .O(x46_y43),
    .I0(x43_y46),
    .I1(1'b0),
    .I2(x44_y42),
    .I3(x43_y48)
);

(* keep, dont_touch *)
(* LOC = "X47/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110010111100)
) lut_47_43 (
    .O(x47_y43),
    .I0(x44_y41),
    .I1(x45_y43),
    .I2(1'b0),
    .I3(x44_y44)
);

(* keep, dont_touch *)
(* LOC = "X48/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101100000110)
) lut_48_43 (
    .O(x48_y43),
    .I0(x46_y47),
    .I1(x46_y47),
    .I2(x46_y38),
    .I3(x45_y48)
);

(* keep, dont_touch *)
(* LOC = "X49/Y43" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101011001110)
) lut_49_43 (
    .O(x49_y43),
    .I0(1'b0),
    .I1(x47_y38),
    .I2(x47_y44),
    .I3(x47_y44)
);

(* keep, dont_touch *)
(* LOC = "X0/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010011010011)
) lut_0_44 (
    .O(x0_y44),
    .I0(in9),
    .I1(in5),
    .I2(1'b0),
    .I3(in0)
);

(* keep, dont_touch *)
(* LOC = "X1/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011001011101)
) lut_1_44 (
    .O(x1_y44),
    .I0(in6),
    .I1(in6),
    .I2(in5),
    .I3(in5)
);

(* keep, dont_touch *)
(* LOC = "X2/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101010001000)
) lut_2_44 (
    .O(x2_y44),
    .I0(in9),
    .I1(1'b0),
    .I2(1'b0),
    .I3(in2)
);

(* keep, dont_touch *)
(* LOC = "X3/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010010001011)
) lut_3_44 (
    .O(x3_y44),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x1_y40),
    .I3(x1_y39)
);

(* keep, dont_touch *)
(* LOC = "X4/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001011010101)
) lut_4_44 (
    .O(x4_y44),
    .I0(1'b0),
    .I1(x1_y49),
    .I2(x1_y44),
    .I3(x1_y40)
);

(* keep, dont_touch *)
(* LOC = "X5/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101111101111110)
) lut_5_44 (
    .O(x5_y44),
    .I0(x3_y39),
    .I1(x2_y47),
    .I2(x3_y44),
    .I3(x2_y49)
);

(* keep, dont_touch *)
(* LOC = "X6/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100000100001)
) lut_6_44 (
    .O(x6_y44),
    .I0(1'b0),
    .I1(x4_y40),
    .I2(x4_y40),
    .I3(x4_y46)
);

(* keep, dont_touch *)
(* LOC = "X7/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111111001110)
) lut_7_44 (
    .O(x7_y44),
    .I0(x5_y43),
    .I1(x4_y42),
    .I2(1'b0),
    .I3(x5_y39)
);

(* keep, dont_touch *)
(* LOC = "X8/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000000010100)
) lut_8_44 (
    .O(x8_y44),
    .I0(x6_y47),
    .I1(x5_y45),
    .I2(x5_y44),
    .I3(x6_y47)
);

(* keep, dont_touch *)
(* LOC = "X9/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000000001100)
) lut_9_44 (
    .O(x9_y44),
    .I0(1'b0),
    .I1(x6_y43),
    .I2(x5_y44),
    .I3(x6_y47)
);

(* keep, dont_touch *)
(* LOC = "X10/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011101000111)
) lut_10_44 (
    .O(x10_y44),
    .I0(x8_y46),
    .I1(x7_y48),
    .I2(x8_y42),
    .I3(x8_y47)
);

(* keep, dont_touch *)
(* LOC = "X11/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111010110111)
) lut_11_44 (
    .O(x11_y44),
    .I0(x9_y40),
    .I1(x8_y39),
    .I2(x8_y39),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X12/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000001110011)
) lut_12_44 (
    .O(x12_y44),
    .I0(1'b0),
    .I1(x9_y43),
    .I2(x9_y48),
    .I3(x9_y42)
);

(* keep, dont_touch *)
(* LOC = "X13/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111001101010)
) lut_13_44 (
    .O(x13_y44),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x10_y49),
    .I3(x10_y41)
);

(* keep, dont_touch *)
(* LOC = "X14/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011000001111011)
) lut_14_44 (
    .O(x14_y44),
    .I0(1'b0),
    .I1(x12_y49),
    .I2(x11_y45),
    .I3(x12_y45)
);

(* keep, dont_touch *)
(* LOC = "X15/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001110011011101)
) lut_15_44 (
    .O(x15_y44),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x13_y48),
    .I3(x12_y41)
);

(* keep, dont_touch *)
(* LOC = "X16/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100011111001)
) lut_16_44 (
    .O(x16_y44),
    .I0(1'b0),
    .I1(x14_y46),
    .I2(x13_y48),
    .I3(x14_y43)
);

(* keep, dont_touch *)
(* LOC = "X17/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011010111101100)
) lut_17_44 (
    .O(x17_y44),
    .I0(x14_y39),
    .I1(x14_y39),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X18/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111011010000)
) lut_18_44 (
    .O(x18_y44),
    .I0(1'b0),
    .I1(x15_y41),
    .I2(x15_y40),
    .I3(x16_y44)
);

(* keep, dont_touch *)
(* LOC = "X19/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011011110000)
) lut_19_44 (
    .O(x19_y44),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x17_y44)
);

(* keep, dont_touch *)
(* LOC = "X20/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001010001000001)
) lut_20_44 (
    .O(x20_y44),
    .I0(x18_y40),
    .I1(x17_y45),
    .I2(x18_y46),
    .I3(x17_y39)
);

(* keep, dont_touch *)
(* LOC = "X21/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000100100000)
) lut_21_44 (
    .O(x21_y44),
    .I0(x18_y49),
    .I1(x18_y47),
    .I2(x18_y39),
    .I3(x18_y41)
);

(* keep, dont_touch *)
(* LOC = "X22/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101111001001)
) lut_22_44 (
    .O(x22_y44),
    .I0(x20_y49),
    .I1(x20_y45),
    .I2(x19_y44),
    .I3(x20_y39)
);

(* keep, dont_touch *)
(* LOC = "X23/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101101001101)
) lut_23_44 (
    .O(x23_y44),
    .I0(x20_y49),
    .I1(x21_y48),
    .I2(1'b0),
    .I3(x21_y41)
);

(* keep, dont_touch *)
(* LOC = "X24/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110110110111)
) lut_24_44 (
    .O(x24_y44),
    .I0(x21_y43),
    .I1(x21_y43),
    .I2(x22_y42),
    .I3(x22_y47)
);

(* keep, dont_touch *)
(* LOC = "X25/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100000000111)
) lut_25_44 (
    .O(x25_y44),
    .I0(x22_y45),
    .I1(x22_y49),
    .I2(x23_y42),
    .I3(x22_y49)
);

(* keep, dont_touch *)
(* LOC = "X26/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110000100010)
) lut_26_44 (
    .O(x26_y44),
    .I0(x23_y47),
    .I1(x24_y43),
    .I2(1'b0),
    .I3(x24_y42)
);

(* keep, dont_touch *)
(* LOC = "X27/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100001010011)
) lut_27_44 (
    .O(x27_y44),
    .I0(x24_y45),
    .I1(1'b0),
    .I2(x24_y44),
    .I3(x25_y49)
);

(* keep, dont_touch *)
(* LOC = "X28/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010101110000)
) lut_28_44 (
    .O(x28_y44),
    .I0(x26_y45),
    .I1(1'b0),
    .I2(x25_y39),
    .I3(x26_y49)
);

(* keep, dont_touch *)
(* LOC = "X29/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101010111010)
) lut_29_44 (
    .O(x29_y44),
    .I0(x27_y44),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X30/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010000011010)
) lut_30_44 (
    .O(x30_y44),
    .I0(x28_y39),
    .I1(x27_y46),
    .I2(x27_y42),
    .I3(x27_y48)
);

(* keep, dont_touch *)
(* LOC = "X31/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111000101000011)
) lut_31_44 (
    .O(x31_y44),
    .I0(x28_y42),
    .I1(x29_y41),
    .I2(x29_y48),
    .I3(x28_y47)
);

(* keep, dont_touch *)
(* LOC = "X32/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111111001000)
) lut_32_44 (
    .O(x32_y44),
    .I0(x30_y44),
    .I1(1'b0),
    .I2(x29_y44),
    .I3(x29_y44)
);

(* keep, dont_touch *)
(* LOC = "X33/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111100110101)
) lut_33_44 (
    .O(x33_y44),
    .I0(x31_y48),
    .I1(x30_y41),
    .I2(x31_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X34/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010111001011)
) lut_34_44 (
    .O(x34_y44),
    .I0(x32_y41),
    .I1(x32_y43),
    .I2(x31_y41),
    .I3(x32_y44)
);

(* keep, dont_touch *)
(* LOC = "X35/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001111110001)
) lut_35_44 (
    .O(x35_y44),
    .I0(1'b0),
    .I1(x33_y41),
    .I2(x32_y40),
    .I3(x32_y42)
);

(* keep, dont_touch *)
(* LOC = "X36/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000110000001)
) lut_36_44 (
    .O(x36_y44),
    .I0(x34_y43),
    .I1(x34_y46),
    .I2(x33_y48),
    .I3(x34_y44)
);

(* keep, dont_touch *)
(* LOC = "X37/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111110001111)
) lut_37_44 (
    .O(x37_y44),
    .I0(x35_y47),
    .I1(x35_y41),
    .I2(x34_y49),
    .I3(x35_y47)
);

(* keep, dont_touch *)
(* LOC = "X38/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101110110010)
) lut_38_44 (
    .O(x38_y44),
    .I0(x35_y45),
    .I1(x36_y47),
    .I2(x35_y48),
    .I3(x35_y39)
);

(* keep, dont_touch *)
(* LOC = "X39/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100011101100111)
) lut_39_44 (
    .O(x39_y44),
    .I0(x36_y43),
    .I1(1'b0),
    .I2(x37_y42),
    .I3(x36_y45)
);

(* keep, dont_touch *)
(* LOC = "X40/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110001010001)
) lut_40_44 (
    .O(x40_y44),
    .I0(x37_y46),
    .I1(x37_y48),
    .I2(x38_y43),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X41/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101110110111)
) lut_41_44 (
    .O(x41_y44),
    .I0(x38_y44),
    .I1(x38_y40),
    .I2(x38_y49),
    .I3(x38_y43)
);

(* keep, dont_touch *)
(* LOC = "X42/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010100100011)
) lut_42_44 (
    .O(x42_y44),
    .I0(x39_y45),
    .I1(x39_y39),
    .I2(x40_y39),
    .I3(x39_y48)
);

(* keep, dont_touch *)
(* LOC = "X43/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001010000000)
) lut_43_44 (
    .O(x43_y44),
    .I0(x41_y43),
    .I1(1'b0),
    .I2(x40_y46),
    .I3(x41_y40)
);

(* keep, dont_touch *)
(* LOC = "X44/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100010110001)
) lut_44_44 (
    .O(x44_y44),
    .I0(x41_y45),
    .I1(1'b0),
    .I2(x41_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X45/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101010010100)
) lut_45_44 (
    .O(x45_y44),
    .I0(x43_y42),
    .I1(x42_y46),
    .I2(x42_y41),
    .I3(x42_y40)
);

(* keep, dont_touch *)
(* LOC = "X46/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001000111010111)
) lut_46_44 (
    .O(x46_y44),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x43_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X47/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110111000110)
) lut_47_44 (
    .O(x47_y44),
    .I0(1'b0),
    .I1(x45_y47),
    .I2(x44_y49),
    .I3(x44_y49)
);

(* keep, dont_touch *)
(* LOC = "X48/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101101011111)
) lut_48_44 (
    .O(x48_y44),
    .I0(x45_y47),
    .I1(x45_y40),
    .I2(x46_y43),
    .I3(x46_y41)
);

(* keep, dont_touch *)
(* LOC = "X49/Y44" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100100110000)
) lut_49_44 (
    .O(x49_y44),
    .I0(x46_y40),
    .I1(x47_y46),
    .I2(1'b0),
    .I3(x46_y48)
);

(* keep, dont_touch *)
(* LOC = "X0/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111000010100)
) lut_0_45 (
    .O(x0_y45),
    .I0(in5),
    .I1(in9),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X1/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010011011101)
) lut_1_45 (
    .O(x1_y45),
    .I0(in4),
    .I1(in7),
    .I2(1'b0),
    .I3(in1)
);

(* keep, dont_touch *)
(* LOC = "X2/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000100010000)
) lut_2_45 (
    .O(x2_y45),
    .I0(1'b0),
    .I1(in5),
    .I2(1'b0),
    .I3(in6)
);

(* keep, dont_touch *)
(* LOC = "X3/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111101110101)
) lut_3_45 (
    .O(x3_y45),
    .I0(in9),
    .I1(1'b0),
    .I2(in9),
    .I3(x1_y45)
);

(* keep, dont_touch *)
(* LOC = "X4/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010011111001)
) lut_4_45 (
    .O(x4_y45),
    .I0(x2_y46),
    .I1(x2_y43),
    .I2(x2_y43),
    .I3(x2_y42)
);

(* keep, dont_touch *)
(* LOC = "X5/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101001011001)
) lut_5_45 (
    .O(x5_y45),
    .I0(x3_y42),
    .I1(x2_y44),
    .I2(1'b0),
    .I3(x2_y49)
);

(* keep, dont_touch *)
(* LOC = "X6/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101110100100)
) lut_6_45 (
    .O(x6_y45),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x3_y40),
    .I3(x4_y47)
);

(* keep, dont_touch *)
(* LOC = "X7/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001001011010111)
) lut_7_45 (
    .O(x7_y45),
    .I0(x5_y49),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X8/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000111111000)
) lut_8_45 (
    .O(x8_y45),
    .I0(x6_y45),
    .I1(x5_y48),
    .I2(x6_y46),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X9/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101111000011)
) lut_9_45 (
    .O(x9_y45),
    .I0(1'b0),
    .I1(x6_y49),
    .I2(x6_y46),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X10/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001011001001)
) lut_10_45 (
    .O(x10_y45),
    .I0(x8_y44),
    .I1(x7_y40),
    .I2(x7_y49),
    .I3(x7_y47)
);

(* keep, dont_touch *)
(* LOC = "X11/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111000001010)
) lut_11_45 (
    .O(x11_y45),
    .I0(1'b0),
    .I1(x9_y40),
    .I2(x9_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X12/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001000010101010)
) lut_12_45 (
    .O(x12_y45),
    .I0(1'b0),
    .I1(x9_y41),
    .I2(1'b0),
    .I3(x9_y40)
);

(* keep, dont_touch *)
(* LOC = "X13/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000001010001)
) lut_13_45 (
    .O(x13_y45),
    .I0(x10_y49),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X14/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110101010111)
) lut_14_45 (
    .O(x14_y45),
    .I0(1'b0),
    .I1(x12_y40),
    .I2(1'b0),
    .I3(x12_y43)
);

(* keep, dont_touch *)
(* LOC = "X15/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100101111001)
) lut_15_45 (
    .O(x15_y45),
    .I0(1'b0),
    .I1(x13_y40),
    .I2(x13_y49),
    .I3(x12_y46)
);

(* keep, dont_touch *)
(* LOC = "X16/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000011010000)
) lut_16_45 (
    .O(x16_y45),
    .I0(x13_y44),
    .I1(1'b0),
    .I2(x14_y45),
    .I3(x13_y46)
);

(* keep, dont_touch *)
(* LOC = "X17/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000010010000010)
) lut_17_45 (
    .O(x17_y45),
    .I0(x14_y48),
    .I1(x15_y45),
    .I2(x14_y47),
    .I3(x15_y45)
);

(* keep, dont_touch *)
(* LOC = "X18/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001100010010)
) lut_18_45 (
    .O(x18_y45),
    .I0(x16_y42),
    .I1(x16_y47),
    .I2(x15_y48),
    .I3(x16_y48)
);

(* keep, dont_touch *)
(* LOC = "X19/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001100100111)
) lut_19_45 (
    .O(x19_y45),
    .I0(x16_y41),
    .I1(x16_y41),
    .I2(1'b0),
    .I3(x16_y41)
);

(* keep, dont_touch *)
(* LOC = "X20/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110010100010100)
) lut_20_45 (
    .O(x20_y45),
    .I0(x18_y41),
    .I1(x18_y40),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X21/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010001110011)
) lut_21_45 (
    .O(x21_y45),
    .I0(x18_y48),
    .I1(x18_y47),
    .I2(1'b0),
    .I3(x18_y43)
);

(* keep, dont_touch *)
(* LOC = "X22/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000001110000)
) lut_22_45 (
    .O(x22_y45),
    .I0(1'b0),
    .I1(x20_y42),
    .I2(x20_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X23/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001011001100)
) lut_23_45 (
    .O(x23_y45),
    .I0(x21_y44),
    .I1(x20_y41),
    .I2(x21_y46),
    .I3(x20_y46)
);

(* keep, dont_touch *)
(* LOC = "X24/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111010000100)
) lut_24_45 (
    .O(x24_y45),
    .I0(x22_y46),
    .I1(x22_y43),
    .I2(1'b0),
    .I3(x22_y43)
);

(* keep, dont_touch *)
(* LOC = "X25/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110100000111)
) lut_25_45 (
    .O(x25_y45),
    .I0(x23_y48),
    .I1(x22_y49),
    .I2(x23_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X26/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001100100000101)
) lut_26_45 (
    .O(x26_y45),
    .I0(1'b0),
    .I1(x24_y48),
    .I2(x23_y41),
    .I3(x24_y41)
);

(* keep, dont_touch *)
(* LOC = "X27/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110101100101)
) lut_27_45 (
    .O(x27_y45),
    .I0(x24_y44),
    .I1(x25_y43),
    .I2(x25_y44),
    .I3(x24_y45)
);

(* keep, dont_touch *)
(* LOC = "X28/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111111100010)
) lut_28_45 (
    .O(x28_y45),
    .I0(x26_y44),
    .I1(x26_y41),
    .I2(x25_y43),
    .I3(x25_y47)
);

(* keep, dont_touch *)
(* LOC = "X29/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101000101101)
) lut_29_45 (
    .O(x29_y45),
    .I0(x26_y48),
    .I1(1'b0),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X30/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101000101101)
) lut_30_45 (
    .O(x30_y45),
    .I0(1'b0),
    .I1(x28_y49),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X31/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101110010101)
) lut_31_45 (
    .O(x31_y45),
    .I0(x28_y49),
    .I1(1'b0),
    .I2(x28_y40),
    .I3(x28_y42)
);

(* keep, dont_touch *)
(* LOC = "X32/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110000001000)
) lut_32_45 (
    .O(x32_y45),
    .I0(x29_y43),
    .I1(x30_y42),
    .I2(x29_y49),
    .I3(x30_y40)
);

(* keep, dont_touch *)
(* LOC = "X33/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101100000000)
) lut_33_45 (
    .O(x33_y45),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x30_y41),
    .I3(x30_y48)
);

(* keep, dont_touch *)
(* LOC = "X34/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101101101011)
) lut_34_45 (
    .O(x34_y45),
    .I0(x32_y40),
    .I1(x31_y49),
    .I2(x31_y49),
    .I3(x31_y45)
);

(* keep, dont_touch *)
(* LOC = "X35/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010011001010)
) lut_35_45 (
    .O(x35_y45),
    .I0(1'b0),
    .I1(x33_y45),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X36/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101101000010)
) lut_36_45 (
    .O(x36_y45),
    .I0(x34_y47),
    .I1(x33_y41),
    .I2(x34_y48),
    .I3(x33_y43)
);

(* keep, dont_touch *)
(* LOC = "X37/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011101010101001)
) lut_37_45 (
    .O(x37_y45),
    .I0(x34_y49),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x35_y42)
);

(* keep, dont_touch *)
(* LOC = "X38/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100100111011)
) lut_38_45 (
    .O(x38_y45),
    .I0(x35_y47),
    .I1(x35_y46),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X39/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110111001100)
) lut_39_45 (
    .O(x39_y45),
    .I0(x36_y45),
    .I1(x37_y44),
    .I2(x36_y48),
    .I3(x37_y47)
);

(* keep, dont_touch *)
(* LOC = "X40/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101111101010)
) lut_40_45 (
    .O(x40_y45),
    .I0(x38_y42),
    .I1(x38_y41),
    .I2(x37_y49),
    .I3(x38_y43)
);

(* keep, dont_touch *)
(* LOC = "X41/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111101100011)
) lut_41_45 (
    .O(x41_y45),
    .I0(x39_y47),
    .I1(x39_y41),
    .I2(x39_y42),
    .I3(x38_y49)
);

(* keep, dont_touch *)
(* LOC = "X42/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110001001011)
) lut_42_45 (
    .O(x42_y45),
    .I0(1'b0),
    .I1(x40_y48),
    .I2(x40_y43),
    .I3(x40_y40)
);

(* keep, dont_touch *)
(* LOC = "X43/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111110111001)
) lut_43_45 (
    .O(x43_y45),
    .I0(1'b0),
    .I1(x41_y48),
    .I2(1'b0),
    .I3(x40_y47)
);

(* keep, dont_touch *)
(* LOC = "X44/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101000010111)
) lut_44_45 (
    .O(x44_y45),
    .I0(x42_y40),
    .I1(x41_y43),
    .I2(1'b0),
    .I3(x42_y44)
);

(* keep, dont_touch *)
(* LOC = "X45/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100110010110)
) lut_45_45 (
    .O(x45_y45),
    .I0(x42_y47),
    .I1(x42_y49),
    .I2(x42_y49),
    .I3(x43_y42)
);

(* keep, dont_touch *)
(* LOC = "X46/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111111001110)
) lut_46_45 (
    .O(x46_y45),
    .I0(x43_y45),
    .I1(1'b0),
    .I2(x43_y43),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X47/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001000111000)
) lut_47_45 (
    .O(x47_y45),
    .I0(x45_y47),
    .I1(x45_y49),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X48/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111000010110)
) lut_48_45 (
    .O(x48_y45),
    .I0(x46_y44),
    .I1(x45_y49),
    .I2(x45_y49),
    .I3(x46_y45)
);

(* keep, dont_touch *)
(* LOC = "X49/Y45" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001100010111)
) lut_49_45 (
    .O(x49_y45),
    .I0(x47_y48),
    .I1(1'b0),
    .I2(x46_y49),
    .I3(x47_y44)
);

(* keep, dont_touch *)
(* LOC = "X0/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011100111111)
) lut_0_46 (
    .O(x0_y46),
    .I0(in9),
    .I1(in3),
    .I2(1'b0),
    .I3(in4)
);

(* keep, dont_touch *)
(* LOC = "X1/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111011001001)
) lut_1_46 (
    .O(x1_y46),
    .I0(in9),
    .I1(in3),
    .I2(1'b0),
    .I3(in9)
);

(* keep, dont_touch *)
(* LOC = "X2/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011000111001)
) lut_2_46 (
    .O(x2_y46),
    .I0(in4),
    .I1(in4),
    .I2(in3),
    .I3(in4)
);

(* keep, dont_touch *)
(* LOC = "X3/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101101100000000)
) lut_3_46 (
    .O(x3_y46),
    .I0(in5),
    .I1(in9),
    .I2(in9),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X4/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010110100000)
) lut_4_46 (
    .O(x4_y46),
    .I0(x2_y46),
    .I1(x1_y49),
    .I2(x2_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X5/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011100001101)
) lut_5_46 (
    .O(x5_y46),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x2_y49),
    .I3(x2_y41)
);

(* keep, dont_touch *)
(* LOC = "X6/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000001011000)
) lut_6_46 (
    .O(x6_y46),
    .I0(1'b0),
    .I1(x4_y49),
    .I2(x3_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X7/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000000110011)
) lut_7_46 (
    .O(x7_y46),
    .I0(x4_y41),
    .I1(x4_y47),
    .I2(1'b0),
    .I3(x4_y49)
);

(* keep, dont_touch *)
(* LOC = "X8/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001111000101)
) lut_8_46 (
    .O(x8_y46),
    .I0(x5_y49),
    .I1(1'b0),
    .I2(x6_y49),
    .I3(x6_y41)
);

(* keep, dont_touch *)
(* LOC = "X9/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011110000111)
) lut_9_46 (
    .O(x9_y46),
    .I0(x7_y43),
    .I1(x6_y42),
    .I2(x6_y49),
    .I3(x6_y41)
);

(* keep, dont_touch *)
(* LOC = "X10/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110001001110)
) lut_10_46 (
    .O(x10_y46),
    .I0(x7_y44),
    .I1(1'b0),
    .I2(x8_y47),
    .I3(x8_y45)
);

(* keep, dont_touch *)
(* LOC = "X11/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000110111100)
) lut_11_46 (
    .O(x11_y46),
    .I0(x8_y48),
    .I1(x8_y48),
    .I2(x9_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X12/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101101101011)
) lut_12_46 (
    .O(x12_y46),
    .I0(1'b0),
    .I1(x9_y41),
    .I2(1'b0),
    .I3(x9_y49)
);

(* keep, dont_touch *)
(* LOC = "X13/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100110110110)
) lut_13_46 (
    .O(x13_y46),
    .I0(x10_y46),
    .I1(x10_y49),
    .I2(x10_y43),
    .I3(x10_y46)
);

(* keep, dont_touch *)
(* LOC = "X14/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101000100000)
) lut_14_46 (
    .O(x14_y46),
    .I0(x12_y41),
    .I1(x12_y48),
    .I2(1'b0),
    .I3(x12_y49)
);

(* keep, dont_touch *)
(* LOC = "X15/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110010010001)
) lut_15_46 (
    .O(x15_y46),
    .I0(1'b0),
    .I1(x12_y42),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X16/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110011000001)
) lut_16_46 (
    .O(x16_y46),
    .I0(1'b0),
    .I1(x14_y46),
    .I2(1'b0),
    .I3(x13_y42)
);

(* keep, dont_touch *)
(* LOC = "X17/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011100111111)
) lut_17_46 (
    .O(x17_y46),
    .I0(x15_y42),
    .I1(x14_y49),
    .I2(x14_y41),
    .I3(x14_y43)
);

(* keep, dont_touch *)
(* LOC = "X18/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011110110110)
) lut_18_46 (
    .O(x18_y46),
    .I0(1'b0),
    .I1(x16_y41),
    .I2(1'b0),
    .I3(x16_y41)
);

(* keep, dont_touch *)
(* LOC = "X19/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010011001100)
) lut_19_46 (
    .O(x19_y46),
    .I0(1'b0),
    .I1(x16_y42),
    .I2(x16_y47),
    .I3(x17_y49)
);

(* keep, dont_touch *)
(* LOC = "X20/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110100010101)
) lut_20_46 (
    .O(x20_y46),
    .I0(x17_y42),
    .I1(1'b0),
    .I2(x17_y49),
    .I3(x17_y43)
);

(* keep, dont_touch *)
(* LOC = "X21/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110110100100)
) lut_21_46 (
    .O(x21_y46),
    .I0(x19_y41),
    .I1(1'b0),
    .I2(x19_y49),
    .I3(x18_y49)
);

(* keep, dont_touch *)
(* LOC = "X22/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100000101011)
) lut_22_46 (
    .O(x22_y46),
    .I0(x20_y42),
    .I1(x19_y46),
    .I2(x20_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X23/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010100001100)
) lut_23_46 (
    .O(x23_y46),
    .I0(x21_y42),
    .I1(x21_y49),
    .I2(x21_y43),
    .I3(x20_y42)
);

(* keep, dont_touch *)
(* LOC = "X24/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101100000101)
) lut_24_46 (
    .O(x24_y46),
    .I0(x22_y49),
    .I1(1'b0),
    .I2(x22_y43),
    .I3(x22_y48)
);

(* keep, dont_touch *)
(* LOC = "X25/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010000000001101)
) lut_25_46 (
    .O(x25_y46),
    .I0(x23_y43),
    .I1(1'b0),
    .I2(x23_y43),
    .I3(x22_y49)
);

(* keep, dont_touch *)
(* LOC = "X26/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001010011001)
) lut_26_46 (
    .O(x26_y46),
    .I0(x23_y42),
    .I1(x23_y43),
    .I2(x23_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X27/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100001110000)
) lut_27_46 (
    .O(x27_y46),
    .I0(x24_y41),
    .I1(x25_y47),
    .I2(x24_y45),
    .I3(x25_y41)
);

(* keep, dont_touch *)
(* LOC = "X28/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110011000111100)
) lut_28_46 (
    .O(x28_y46),
    .I0(x25_y45),
    .I1(x25_y44),
    .I2(x26_y43),
    .I3(x26_y49)
);

(* keep, dont_touch *)
(* LOC = "X29/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010111011000)
) lut_29_46 (
    .O(x29_y46),
    .I0(x27_y48),
    .I1(x26_y47),
    .I2(1'b0),
    .I3(x26_y44)
);

(* keep, dont_touch *)
(* LOC = "X30/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110111000001)
) lut_30_46 (
    .O(x30_y46),
    .I0(x27_y49),
    .I1(x27_y48),
    .I2(x28_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X31/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101001011111001)
) lut_31_46 (
    .O(x31_y46),
    .I0(x28_y49),
    .I1(x29_y49),
    .I2(x29_y45),
    .I3(x29_y49)
);

(* keep, dont_touch *)
(* LOC = "X32/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010101110001)
) lut_32_46 (
    .O(x32_y46),
    .I0(1'b0),
    .I1(x30_y43),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X33/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001001101110001)
) lut_33_46 (
    .O(x33_y46),
    .I0(x30_y48),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x31_y43)
);

(* keep, dont_touch *)
(* LOC = "X34/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100000101101101)
) lut_34_46 (
    .O(x34_y46),
    .I0(x32_y49),
    .I1(1'b0),
    .I2(x32_y46),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X35/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111111011000000)
) lut_35_46 (
    .O(x35_y46),
    .I0(x33_y47),
    .I1(x32_y44),
    .I2(x32_y43),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X36/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111101100010)
) lut_36_46 (
    .O(x36_y46),
    .I0(x33_y49),
    .I1(1'b0),
    .I2(x33_y46),
    .I3(x33_y43)
);

(* keep, dont_touch *)
(* LOC = "X37/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111101011001111)
) lut_37_46 (
    .O(x37_y46),
    .I0(x34_y49),
    .I1(x35_y48),
    .I2(1'b0),
    .I3(x35_y46)
);

(* keep, dont_touch *)
(* LOC = "X38/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000001110000111)
) lut_38_46 (
    .O(x38_y46),
    .I0(x35_y49),
    .I1(x36_y43),
    .I2(x36_y45),
    .I3(x36_y42)
);

(* keep, dont_touch *)
(* LOC = "X39/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111100001010011)
) lut_39_46 (
    .O(x39_y46),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x37_y49),
    .I3(x37_y43)
);

(* keep, dont_touch *)
(* LOC = "X40/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100001000000010)
) lut_40_46 (
    .O(x40_y46),
    .I0(x37_y48),
    .I1(x37_y41),
    .I2(x38_y43),
    .I3(x37_y45)
);

(* keep, dont_touch *)
(* LOC = "X41/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011111011111011)
) lut_41_46 (
    .O(x41_y46),
    .I0(x39_y44),
    .I1(1'b0),
    .I2(x39_y49),
    .I3(x38_y41)
);

(* keep, dont_touch *)
(* LOC = "X42/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111011000011)
) lut_42_46 (
    .O(x42_y46),
    .I0(1'b0),
    .I1(x39_y49),
    .I2(x39_y49),
    .I3(x39_y48)
);

(* keep, dont_touch *)
(* LOC = "X43/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111100011010)
) lut_43_46 (
    .O(x43_y46),
    .I0(x40_y49),
    .I1(1'b0),
    .I2(x40_y49),
    .I3(x40_y48)
);

(* keep, dont_touch *)
(* LOC = "X44/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111010011001010)
) lut_44_46 (
    .O(x44_y46),
    .I0(x41_y45),
    .I1(x41_y44),
    .I2(x42_y49),
    .I3(x41_y43)
);

(* keep, dont_touch *)
(* LOC = "X45/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111110110101)
) lut_45_46 (
    .O(x45_y46),
    .I0(x42_y44),
    .I1(x43_y44),
    .I2(x43_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X46/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011101110001)
) lut_46_46 (
    .O(x46_y46),
    .I0(x43_y48),
    .I1(x43_y46),
    .I2(x43_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X47/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011100101011001)
) lut_47_46 (
    .O(x47_y46),
    .I0(x45_y49),
    .I1(x44_y49),
    .I2(x44_y44),
    .I3(x45_y44)
);

(* keep, dont_touch *)
(* LOC = "X48/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100101000001)
) lut_48_46 (
    .O(x48_y46),
    .I0(1'b0),
    .I1(x46_y45),
    .I2(x45_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X49/Y46" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110000110101010)
) lut_49_46 (
    .O(x49_y46),
    .I0(x47_y46),
    .I1(x46_y45),
    .I2(1'b0),
    .I3(x46_y47)
);

(* keep, dont_touch *)
(* LOC = "X0/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110010111001)
) lut_0_47 (
    .O(x0_y47),
    .I0(in2),
    .I1(1'b0),
    .I2(in7),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X1/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100100000110)
) lut_1_47 (
    .O(x1_y47),
    .I0(in9),
    .I1(in8),
    .I2(in8),
    .I3(in2)
);

(* keep, dont_touch *)
(* LOC = "X2/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100101101010)
) lut_2_47 (
    .O(x2_y47),
    .I0(in9),
    .I1(in3),
    .I2(in5),
    .I3(in9)
);

(* keep, dont_touch *)
(* LOC = "X3/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101100100110)
) lut_3_47 (
    .O(x3_y47),
    .I0(in9),
    .I1(x1_y46),
    .I2(x1_y44),
    .I3(in4)
);

(* keep, dont_touch *)
(* LOC = "X4/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111011010101010)
) lut_4_47 (
    .O(x4_y47),
    .I0(x1_y48),
    .I1(x1_y45),
    .I2(x1_y42),
    .I3(x2_y44)
);

(* keep, dont_touch *)
(* LOC = "X5/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001100110000101)
) lut_5_47 (
    .O(x5_y47),
    .I0(x3_y49),
    .I1(x2_y43),
    .I2(1'b0),
    .I3(x2_y49)
);

(* keep, dont_touch *)
(* LOC = "X6/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010010010110)
) lut_6_47 (
    .O(x6_y47),
    .I0(x3_y49),
    .I1(1'b0),
    .I2(x3_y49),
    .I3(x4_y45)
);

(* keep, dont_touch *)
(* LOC = "X7/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010100111000)
) lut_7_47 (
    .O(x7_y47),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x5_y45),
    .I3(x5_y49)
);

(* keep, dont_touch *)
(* LOC = "X8/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101001000011)
) lut_8_47 (
    .O(x8_y47),
    .I0(x6_y49),
    .I1(x5_y49),
    .I2(x6_y49),
    .I3(x6_y49)
);

(* keep, dont_touch *)
(* LOC = "X9/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100100011010)
) lut_9_47 (
    .O(x9_y47),
    .I0(x6_y49),
    .I1(1'b0),
    .I2(x6_y49),
    .I3(x6_y49)
);

(* keep, dont_touch *)
(* LOC = "X10/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111100111000001)
) lut_10_47 (
    .O(x10_y47),
    .I0(x8_y43),
    .I1(x8_y46),
    .I2(x8_y43),
    .I3(x7_y46)
);

(* keep, dont_touch *)
(* LOC = "X11/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000000111001110)
) lut_11_47 (
    .O(x11_y47),
    .I0(x8_y46),
    .I1(x8_y43),
    .I2(x8_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X12/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111001010000)
) lut_12_47 (
    .O(x12_y47),
    .I0(x10_y45),
    .I1(x9_y42),
    .I2(x10_y46),
    .I3(x9_y42)
);

(* keep, dont_touch *)
(* LOC = "X13/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100100111000)
) lut_13_47 (
    .O(x13_y47),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x11_y42),
    .I3(x11_y49)
);

(* keep, dont_touch *)
(* LOC = "X14/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110111001100)
) lut_14_47 (
    .O(x14_y47),
    .I0(1'b0),
    .I1(x11_y46),
    .I2(x11_y44),
    .I3(x11_y49)
);

(* keep, dont_touch *)
(* LOC = "X15/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100111000110)
) lut_15_47 (
    .O(x15_y47),
    .I0(1'b0),
    .I1(x13_y45),
    .I2(x13_y47),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X16/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011100111101110)
) lut_16_47 (
    .O(x16_y47),
    .I0(1'b0),
    .I1(x13_y49),
    .I2(x14_y42),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X17/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011001110100)
) lut_17_47 (
    .O(x17_y47),
    .I0(x15_y49),
    .I1(x15_y49),
    .I2(1'b0),
    .I3(x15_y49)
);

(* keep, dont_touch *)
(* LOC = "X18/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110011000110010)
) lut_18_47 (
    .O(x18_y47),
    .I0(x15_y44),
    .I1(x15_y42),
    .I2(x16_y46),
    .I3(x15_y49)
);

(* keep, dont_touch *)
(* LOC = "X19/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111001001000)
) lut_19_47 (
    .O(x19_y47),
    .I0(x16_y47),
    .I1(x16_y46),
    .I2(x16_y45),
    .I3(x16_y48)
);

(* keep, dont_touch *)
(* LOC = "X20/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110010001011)
) lut_20_47 (
    .O(x20_y47),
    .I0(x17_y49),
    .I1(1'b0),
    .I2(x18_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X21/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110011010111)
) lut_21_47 (
    .O(x21_y47),
    .I0(x18_y49),
    .I1(x19_y49),
    .I2(x18_y49),
    .I3(x19_y49)
);

(* keep, dont_touch *)
(* LOC = "X22/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111001001010)
) lut_22_47 (
    .O(x22_y47),
    .I0(x20_y49),
    .I1(x19_y48),
    .I2(x19_y48),
    .I3(x20_y45)
);

(* keep, dont_touch *)
(* LOC = "X23/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011100001001)
) lut_23_47 (
    .O(x23_y47),
    .I0(x20_y49),
    .I1(x20_y49),
    .I2(x21_y42),
    .I3(x21_y46)
);

(* keep, dont_touch *)
(* LOC = "X24/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111000010101)
) lut_24_47 (
    .O(x24_y47),
    .I0(x21_y46),
    .I1(x21_y49),
    .I2(x22_y47),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X25/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001110110011)
) lut_25_47 (
    .O(x25_y47),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x22_y49),
    .I3(x22_y49)
);

(* keep, dont_touch *)
(* LOC = "X26/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110100010000)
) lut_26_47 (
    .O(x26_y47),
    .I0(x23_y44),
    .I1(x23_y49),
    .I2(x23_y49),
    .I3(x23_y42)
);

(* keep, dont_touch *)
(* LOC = "X27/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001000110011)
) lut_27_47 (
    .O(x27_y47),
    .I0(x24_y42),
    .I1(x24_y43),
    .I2(x25_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X28/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111011101101111)
) lut_28_47 (
    .O(x28_y47),
    .I0(x26_y49),
    .I1(x26_y49),
    .I2(x26_y46),
    .I3(x25_y49)
);

(* keep, dont_touch *)
(* LOC = "X29/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110101110000)
) lut_29_47 (
    .O(x29_y47),
    .I0(x27_y47),
    .I1(x26_y47),
    .I2(1'b0),
    .I3(x27_y49)
);

(* keep, dont_touch *)
(* LOC = "X30/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101100001111111)
) lut_30_47 (
    .O(x30_y47),
    .I0(x28_y49),
    .I1(x28_y47),
    .I2(x28_y43),
    .I3(x27_y47)
);

(* keep, dont_touch *)
(* LOC = "X31/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001010010110001)
) lut_31_47 (
    .O(x31_y47),
    .I0(x29_y49),
    .I1(1'b0),
    .I2(x29_y49),
    .I3(x29_y46)
);

(* keep, dont_touch *)
(* LOC = "X32/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100011011100)
) lut_32_47 (
    .O(x32_y47),
    .I0(1'b0),
    .I1(x30_y42),
    .I2(x29_y42),
    .I3(x30_y44)
);

(* keep, dont_touch *)
(* LOC = "X33/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111000011000)
) lut_33_47 (
    .O(x33_y47),
    .I0(1'b0),
    .I1(x31_y45),
    .I2(x30_y47),
    .I3(x31_y46)
);

(* keep, dont_touch *)
(* LOC = "X34/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111110110011)
) lut_34_47 (
    .O(x34_y47),
    .I0(x32_y49),
    .I1(x31_y44),
    .I2(x32_y42),
    .I3(x32_y46)
);

(* keep, dont_touch *)
(* LOC = "X35/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101110110011)
) lut_35_47 (
    .O(x35_y47),
    .I0(x32_y49),
    .I1(x33_y49),
    .I2(x32_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X36/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010100100000)
) lut_36_47 (
    .O(x36_y47),
    .I0(x34_y49),
    .I1(x33_y48),
    .I2(x33_y42),
    .I3(x33_y49)
);

(* keep, dont_touch *)
(* LOC = "X37/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001000011101)
) lut_37_47 (
    .O(x37_y47),
    .I0(1'b0),
    .I1(x35_y46),
    .I2(x34_y49),
    .I3(x35_y42)
);

(* keep, dont_touch *)
(* LOC = "X38/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010100001110)
) lut_38_47 (
    .O(x38_y47),
    .I0(x36_y49),
    .I1(x35_y46),
    .I2(x35_y49),
    .I3(x35_y49)
);

(* keep, dont_touch *)
(* LOC = "X39/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100011101011)
) lut_39_47 (
    .O(x39_y47),
    .I0(1'b0),
    .I1(x36_y48),
    .I2(x36_y47),
    .I3(x36_y42)
);

(* keep, dont_touch *)
(* LOC = "X40/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000011111000000)
) lut_40_47 (
    .O(x40_y47),
    .I0(x37_y44),
    .I1(x37_y45),
    .I2(x37_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X41/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110010000010)
) lut_41_47 (
    .O(x41_y47),
    .I0(x39_y47),
    .I1(x39_y46),
    .I2(x38_y42),
    .I3(x38_y46)
);

(* keep, dont_touch *)
(* LOC = "X42/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000101110001010)
) lut_42_47 (
    .O(x42_y47),
    .I0(1'b0),
    .I1(x40_y44),
    .I2(x39_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X43/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111101011010)
) lut_43_47 (
    .O(x43_y47),
    .I0(1'b0),
    .I1(x41_y47),
    .I2(1'b0),
    .I3(x41_y48)
);

(* keep, dont_touch *)
(* LOC = "X44/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100001000001000)
) lut_44_47 (
    .O(x44_y47),
    .I0(x42_y42),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x42_y46)
);

(* keep, dont_touch *)
(* LOC = "X45/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011011000000110)
) lut_45_47 (
    .O(x45_y47),
    .I0(x43_y48),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x42_y43)
);

(* keep, dont_touch *)
(* LOC = "X46/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100011010100010)
) lut_46_47 (
    .O(x46_y47),
    .I0(1'b0),
    .I1(x43_y45),
    .I2(x44_y49),
    .I3(x44_y48)
);

(* keep, dont_touch *)
(* LOC = "X47/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010001010110111)
) lut_47_47 (
    .O(x47_y47),
    .I0(x44_y42),
    .I1(1'b0),
    .I2(x45_y49),
    .I3(x45_y43)
);

(* keep, dont_touch *)
(* LOC = "X48/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000111001010)
) lut_48_47 (
    .O(x48_y47),
    .I0(x46_y48),
    .I1(1'b0),
    .I2(x45_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X49/Y47" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100001111001)
) lut_49_47 (
    .O(x49_y47),
    .I0(x47_y46),
    .I1(x47_y45),
    .I2(x46_y47),
    .I3(x46_y49)
);

(* keep, dont_touch *)
(* LOC = "X0/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000111011111111)
) lut_0_48 (
    .O(x0_y48),
    .I0(1'b0),
    .I1(in9),
    .I2(in3),
    .I3(in4)
);

(* keep, dont_touch *)
(* LOC = "X1/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101011110110111)
) lut_1_48 (
    .O(x1_y48),
    .I0(in5),
    .I1(in9),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X2/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001011110011)
) lut_2_48 (
    .O(x2_y48),
    .I0(1'b0),
    .I1(in5),
    .I2(in9),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X3/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100100101010111)
) lut_3_48 (
    .O(x3_y48),
    .I0(in6),
    .I1(in9),
    .I2(1'b0),
    .I3(x1_y49)
);

(* keep, dont_touch *)
(* LOC = "X4/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011000001010)
) lut_4_48 (
    .O(x4_y48),
    .I0(x2_y47),
    .I1(x1_y46),
    .I2(1'b0),
    .I3(x2_y45)
);

(* keep, dont_touch *)
(* LOC = "X5/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110110101010101)
) lut_5_48 (
    .O(x5_y48),
    .I0(x2_y49),
    .I1(x3_y49),
    .I2(1'b0),
    .I3(x2_y49)
);

(* keep, dont_touch *)
(* LOC = "X6/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101001101111101)
) lut_6_48 (
    .O(x6_y48),
    .I0(x4_y43),
    .I1(x3_y49),
    .I2(x3_y43),
    .I3(x4_y49)
);

(* keep, dont_touch *)
(* LOC = "X7/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110110101000)
) lut_7_48 (
    .O(x7_y48),
    .I0(x4_y49),
    .I1(1'b0),
    .I2(x4_y49),
    .I3(x4_y44)
);

(* keep, dont_touch *)
(* LOC = "X8/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000011010000010)
) lut_8_48 (
    .O(x8_y48),
    .I0(x6_y49),
    .I1(x6_y49),
    .I2(x6_y47),
    .I3(x6_y49)
);

(* keep, dont_touch *)
(* LOC = "X9/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000111010001)
) lut_9_48 (
    .O(x9_y48),
    .I0(x6_y47),
    .I1(x7_y49),
    .I2(x6_y47),
    .I3(x6_y49)
);

(* keep, dont_touch *)
(* LOC = "X10/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101100010110)
) lut_10_48 (
    .O(x10_y48),
    .I0(x8_y46),
    .I1(1'b0),
    .I2(x7_y47),
    .I3(x8_y44)
);

(* keep, dont_touch *)
(* LOC = "X11/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101011010010)
) lut_11_48 (
    .O(x11_y48),
    .I0(x9_y48),
    .I1(x9_y47),
    .I2(1'b0),
    .I3(x9_y49)
);

(* keep, dont_touch *)
(* LOC = "X12/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011010101001)
) lut_12_48 (
    .O(x12_y48),
    .I0(x9_y49),
    .I1(x10_y47),
    .I2(x10_y46),
    .I3(x9_y46)
);

(* keep, dont_touch *)
(* LOC = "X13/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110010111111100)
) lut_13_48 (
    .O(x13_y48),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x10_y44),
    .I3(x10_y49)
);

(* keep, dont_touch *)
(* LOC = "X14/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110111100010000)
) lut_14_48 (
    .O(x14_y48),
    .I0(x12_y45),
    .I1(1'b0),
    .I2(x11_y49),
    .I3(x12_y44)
);

(* keep, dont_touch *)
(* LOC = "X15/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111111011001)
) lut_15_48 (
    .O(x15_y48),
    .I0(x13_y49),
    .I1(1'b0),
    .I2(x12_y47),
    .I3(x13_y44)
);

(* keep, dont_touch *)
(* LOC = "X16/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101101111100)
) lut_16_48 (
    .O(x16_y48),
    .I0(x14_y45),
    .I1(x13_y49),
    .I2(x13_y49),
    .I3(x13_y49)
);

(* keep, dont_touch *)
(* LOC = "X17/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110111010000)
) lut_17_48 (
    .O(x17_y48),
    .I0(x14_y49),
    .I1(x14_y47),
    .I2(x15_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X18/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011110000000010)
) lut_18_48 (
    .O(x18_y48),
    .I0(1'b0),
    .I1(x16_y45),
    .I2(x16_y49),
    .I3(x16_y49)
);

(* keep, dont_touch *)
(* LOC = "X19/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101101000101)
) lut_19_48 (
    .O(x19_y48),
    .I0(x16_y44),
    .I1(x17_y48),
    .I2(x17_y49),
    .I3(x17_y46)
);

(* keep, dont_touch *)
(* LOC = "X20/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001101001011)
) lut_20_48 (
    .O(x20_y48),
    .I0(x18_y48),
    .I1(x17_y47),
    .I2(x18_y49),
    .I3(x17_y49)
);

(* keep, dont_touch *)
(* LOC = "X21/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110110101101010)
) lut_21_48 (
    .O(x21_y48),
    .I0(x18_y48),
    .I1(x18_y43),
    .I2(1'b0),
    .I3(x18_y49)
);

(* keep, dont_touch *)
(* LOC = "X22/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011001101111)
) lut_22_48 (
    .O(x22_y48),
    .I0(1'b0),
    .I1(x19_y48),
    .I2(x20_y49),
    .I3(x19_y46)
);

(* keep, dont_touch *)
(* LOC = "X23/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010010011011001)
) lut_23_48 (
    .O(x23_y48),
    .I0(x20_y49),
    .I1(x20_y46),
    .I2(x20_y49),
    .I3(x20_y49)
);

(* keep, dont_touch *)
(* LOC = "X24/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110111110010010)
) lut_24_48 (
    .O(x24_y48),
    .I0(x21_y49),
    .I1(x21_y49),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X25/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000100000010011)
) lut_25_48 (
    .O(x25_y48),
    .I0(x23_y46),
    .I1(x22_y49),
    .I2(x22_y46),
    .I3(x23_y47)
);

(* keep, dont_touch *)
(* LOC = "X26/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001011001110111)
) lut_26_48 (
    .O(x26_y48),
    .I0(x23_y49),
    .I1(x23_y49),
    .I2(x24_y47),
    .I3(x23_y44)
);

(* keep, dont_touch *)
(* LOC = "X27/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100110101110)
) lut_27_48 (
    .O(x27_y48),
    .I0(x24_y48),
    .I1(x25_y45),
    .I2(1'b0),
    .I3(x25_y43)
);

(* keep, dont_touch *)
(* LOC = "X28/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111110111101)
) lut_28_48 (
    .O(x28_y48),
    .I0(x26_y43),
    .I1(x25_y49),
    .I2(x25_y47),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X29/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100111110011010)
) lut_29_48 (
    .O(x29_y48),
    .I0(x26_y45),
    .I1(x27_y49),
    .I2(x27_y43),
    .I3(x26_y47)
);

(* keep, dont_touch *)
(* LOC = "X30/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110101110011001)
) lut_30_48 (
    .O(x30_y48),
    .I0(1'b0),
    .I1(x28_y49),
    .I2(x27_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X31/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101000100000010)
) lut_31_48 (
    .O(x31_y48),
    .I0(x28_y46),
    .I1(x29_y46),
    .I2(1'b0),
    .I3(x28_y47)
);

(* keep, dont_touch *)
(* LOC = "X32/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000010000100010)
) lut_32_48 (
    .O(x32_y48),
    .I0(x30_y49),
    .I1(1'b0),
    .I2(x30_y49),
    .I3(x30_y44)
);

(* keep, dont_touch *)
(* LOC = "X33/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010001000001110)
) lut_33_48 (
    .O(x33_y48),
    .I0(x31_y45),
    .I1(x30_y49),
    .I2(x31_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X34/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001000111110)
) lut_34_48 (
    .O(x34_y48),
    .I0(x31_y46),
    .I1(x32_y48),
    .I2(x32_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X35/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101101001000011)
) lut_35_48 (
    .O(x35_y48),
    .I0(x33_y49),
    .I1(1'b0),
    .I2(x32_y44),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X36/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001101001101)
) lut_36_48 (
    .O(x36_y48),
    .I0(x33_y49),
    .I1(x33_y46),
    .I2(x34_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X37/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101011000011)
) lut_37_48 (
    .O(x37_y48),
    .I0(x34_y44),
    .I1(x35_y43),
    .I2(x34_y49),
    .I3(x34_y43)
);

(* keep, dont_touch *)
(* LOC = "X38/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101010100111)
) lut_38_48 (
    .O(x38_y48),
    .I0(x36_y49),
    .I1(x35_y49),
    .I2(x36_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X39/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0000110001101101)
) lut_39_48 (
    .O(x39_y48),
    .I0(x37_y43),
    .I1(x36_y47),
    .I2(x37_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X40/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010111110101100)
) lut_40_48 (
    .O(x40_y48),
    .I0(x38_y45),
    .I1(x37_y45),
    .I2(x38_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X41/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101101110110)
) lut_41_48 (
    .O(x41_y48),
    .I0(x38_y45),
    .I1(x39_y49),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X42/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111001100001110)
) lut_42_48 (
    .O(x42_y48),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x39_y47),
    .I3(x40_y49)
);

(* keep, dont_touch *)
(* LOC = "X43/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000110111100001)
) lut_43_48 (
    .O(x43_y48),
    .I0(x41_y43),
    .I1(1'b0),
    .I2(x40_y49),
    .I3(x41_y44)
);

(* keep, dont_touch *)
(* LOC = "X44/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101111011100000)
) lut_44_48 (
    .O(x44_y48),
    .I0(1'b0),
    .I1(x42_y49),
    .I2(1'b0),
    .I3(x42_y49)
);

(* keep, dont_touch *)
(* LOC = "X45/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101001001011)
) lut_45_48 (
    .O(x45_y48),
    .I0(x43_y48),
    .I1(x43_y48),
    .I2(1'b0),
    .I3(x43_y49)
);

(* keep, dont_touch *)
(* LOC = "X46/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010110010010011)
) lut_46_48 (
    .O(x46_y48),
    .I0(1'b0),
    .I1(x44_y44),
    .I2(x43_y49),
    .I3(x44_y45)
);

(* keep, dont_touch *)
(* LOC = "X47/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100010010100101)
) lut_47_48 (
    .O(x47_y48),
    .I0(1'b0),
    .I1(1'b0),
    .I2(x45_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X48/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101110111000000)
) lut_48_48 (
    .O(x48_y48),
    .I0(x46_y49),
    .I1(x45_y46),
    .I2(x45_y48),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X49/Y48" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111010111011111)
) lut_49_48 (
    .O(x49_y48),
    .I0(1'b0),
    .I1(x46_y49),
    .I2(x46_y46),
    .I3(x47_y49)
);

(* keep, dont_touch *)
(* LOC = "X0/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011110011100100)
) lut_0_49 (
    .O(x0_y49),
    .I0(in5),
    .I1(1'b0),
    .I2(in9),
    .I3(in9)
);

(* keep, dont_touch *)
(* LOC = "X1/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100000100000111)
) lut_1_49 (
    .O(x1_y49),
    .I0(in9),
    .I1(1'b0),
    .I2(in9),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X2/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011010101101011)
) lut_2_49 (
    .O(x2_y49),
    .I0(1'b0),
    .I1(in7),
    .I2(1'b0),
    .I3(in4)
);

(* keep, dont_touch *)
(* LOC = "X3/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000100001101011)
) lut_3_49 (
    .O(x3_y49),
    .I0(in5),
    .I1(in8),
    .I2(1'b0),
    .I3(x1_y49)
);

(* keep, dont_touch *)
(* LOC = "X4/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100100100101)
) lut_4_49 (
    .O(x4_y49),
    .I0(x2_y48),
    .I1(x2_y44),
    .I2(x2_y45),
    .I3(x2_y49)
);

(* keep, dont_touch *)
(* LOC = "X5/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000111110111100)
) lut_5_49 (
    .O(x5_y49),
    .I0(x3_y47),
    .I1(x2_y44),
    .I2(1'b0),
    .I3(x2_y45)
);

(* keep, dont_touch *)
(* LOC = "X6/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010110000010111)
) lut_6_49 (
    .O(x6_y49),
    .I0(x4_y49),
    .I1(x4_y47),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X7/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010100001101)
) lut_7_49 (
    .O(x7_y49),
    .I0(x5_y49),
    .I1(x5_y45),
    .I2(x4_y49),
    .I3(x4_y44)
);

(* keep, dont_touch *)
(* LOC = "X8/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001101110011001)
) lut_8_49 (
    .O(x8_y49),
    .I0(x6_y48),
    .I1(x6_y49),
    .I2(x5_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X9/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1100101011010101)
) lut_9_49 (
    .O(x9_y49),
    .I0(x6_y48),
    .I1(x7_y49),
    .I2(x5_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X10/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100010110000000)
) lut_10_49 (
    .O(x10_y49),
    .I0(x7_y48),
    .I1(x8_y49),
    .I2(x7_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X11/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111000101000100)
) lut_11_49 (
    .O(x11_y49),
    .I0(1'b0),
    .I1(x9_y49),
    .I2(1'b0),
    .I3(x9_y49)
);

(* keep, dont_touch *)
(* LOC = "X12/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010101100101111)
) lut_12_49 (
    .O(x12_y49),
    .I0(x9_y48),
    .I1(x9_y49),
    .I2(x9_y44),
    .I3(x10_y49)
);

(* keep, dont_touch *)
(* LOC = "X13/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011000000011100)
) lut_13_49 (
    .O(x13_y49),
    .I0(1'b0),
    .I1(x10_y49),
    .I2(1'b0),
    .I3(x11_y49)
);

(* keep, dont_touch *)
(* LOC = "X14/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100100010111110)
) lut_14_49 (
    .O(x14_y49),
    .I0(x11_y49),
    .I1(x12_y49),
    .I2(x12_y49),
    .I3(x12_y49)
);

(* keep, dont_touch *)
(* LOC = "X15/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001101011010011)
) lut_15_49 (
    .O(x15_y49),
    .I0(x12_y49),
    .I1(x13_y49),
    .I2(x13_y49),
    .I3(x13_y49)
);

(* keep, dont_touch *)
(* LOC = "X16/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000001111101111)
) lut_16_49 (
    .O(x16_y49),
    .I0(x14_y45),
    .I1(x14_y44),
    .I2(x14_y46),
    .I3(x14_y48)
);

(* keep, dont_touch *)
(* LOC = "X17/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111010111110)
) lut_17_49 (
    .O(x17_y49),
    .I0(x15_y49),
    .I1(x15_y49),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X18/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1001011000100101)
) lut_18_49 (
    .O(x18_y49),
    .I0(1'b0),
    .I1(x15_y49),
    .I2(x15_y49),
    .I3(x16_y49)
);

(* keep, dont_touch *)
(* LOC = "X19/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001011101110)
) lut_19_49 (
    .O(x19_y49),
    .I0(x17_y44),
    .I1(x16_y45),
    .I2(x16_y48),
    .I3(x16_y48)
);

(* keep, dont_touch *)
(* LOC = "X20/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110011010111)
) lut_20_49 (
    .O(x20_y49),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x18_y49)
);

(* keep, dont_touch *)
(* LOC = "X21/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011011010000010)
) lut_21_49 (
    .O(x21_y49),
    .I0(1'b0),
    .I1(1'b0),
    .I2(1'b0),
    .I3(x19_y48)
);

(* keep, dont_touch *)
(* LOC = "X22/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100001101011)
) lut_22_49 (
    .O(x22_y49),
    .I0(x20_y49),
    .I1(x20_y44),
    .I2(x20_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X23/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110101001010101)
) lut_23_49 (
    .O(x23_y49),
    .I0(x21_y45),
    .I1(x20_y49),
    .I2(x21_y49),
    .I3(x21_y46)
);

(* keep, dont_touch *)
(* LOC = "X24/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1110100111111100)
) lut_24_49 (
    .O(x24_y49),
    .I0(x22_y49),
    .I1(x22_y49),
    .I2(x22_y45),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X25/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111111110011101)
) lut_25_49 (
    .O(x25_y49),
    .I0(x23_y49),
    .I1(x22_y48),
    .I2(x22_y48),
    .I3(x22_y46)
);

(* keep, dont_touch *)
(* LOC = "X26/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b0101100101010110)
) lut_26_49 (
    .O(x26_y49),
    .I0(x23_y49),
    .I1(x23_y49),
    .I2(1'b0),
    .I3(x23_y49)
);

(* keep, dont_touch *)
(* LOC = "X27/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101011001110111)
) lut_27_49 (
    .O(x27_y49),
    .I0(1'b0),
    .I1(x25_y49),
    .I2(1'b0),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X28/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010010101101010)
) lut_28_49 (
    .O(x28_y49),
    .I0(x26_y49),
    .I1(x25_y46),
    .I2(x25_y49),
    .I3(x25_y49)
);

(* keep, dont_touch *)
(* LOC = "X29/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100101111100011)
) lut_29_49 (
    .O(x29_y49),
    .I0(x27_y46),
    .I1(x26_y49),
    .I2(x26_y44),
    .I3(x27_y49)
);

(* keep, dont_touch *)
(* LOC = "X30/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011101100011001)
) lut_30_49 (
    .O(x30_y49),
    .I0(x28_y44),
    .I1(1'b0),
    .I2(x28_y45),
    .I3(x27_y49)
);

(* keep, dont_touch *)
(* LOC = "X31/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011001011101011)
) lut_31_49 (
    .O(x31_y49),
    .I0(x28_y49),
    .I1(1'b0),
    .I2(x28_y49),
    .I3(x29_y46)
);

(* keep, dont_touch *)
(* LOC = "X32/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b0100110000111001)
) lut_32_49 (
    .O(x32_y49),
    .I0(x30_y49),
    .I1(x29_y49),
    .I2(x29_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X33/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1101010111100010)
) lut_33_49 (
    .O(x33_y49),
    .I0(x30_y47),
    .I1(1'b0),
    .I2(x30_y46),
    .I3(x31_y45)
);

(* keep, dont_touch *)
(* LOC = "X34/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111001011011111)
) lut_34_49 (
    .O(x34_y49),
    .I0(1'b0),
    .I1(x31_y49),
    .I2(1'b0),
    .I3(x32_y44)
);

(* keep, dont_touch *)
(* LOC = "X35/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010000110101011)
) lut_35_49 (
    .O(x35_y49),
    .I0(1'b0),
    .I1(x33_y45),
    .I2(x32_y46),
    .I3(x33_y49)
);

(* keep, dont_touch *)
(* LOC = "X36/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010100001100011)
) lut_36_49 (
    .O(x36_y49),
    .I0(x33_y49),
    .I1(1'b0),
    .I2(x33_y49),
    .I3(x33_y49)
);

(* keep, dont_touch *)
(* LOC = "X37/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b0011001111001000)
) lut_37_49 (
    .O(x37_y49),
    .I0(x34_y45),
    .I1(x34_y47),
    .I2(x35_y48),
    .I3(x35_y47)
);

(* keep, dont_touch *)
(* LOC = "X38/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b0110100110000100)
) lut_38_49 (
    .O(x38_y49),
    .I0(x35_y47),
    .I1(x35_y49),
    .I2(1'b0),
    .I3(x35_y49)
);

(* keep, dont_touch *)
(* LOC = "X39/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000000000011)
) lut_39_49 (
    .O(x39_y49),
    .I0(x36_y49),
    .I1(x37_y49),
    .I2(x37_y46),
    .I3(x37_y49)
);

(* keep, dont_touch *)
(* LOC = "X40/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b0001111011100100)
) lut_40_49 (
    .O(x40_y49),
    .I0(1'b0),
    .I1(x38_y45),
    .I2(x37_y47),
    .I3(x38_y49)
);

(* keep, dont_touch *)
(* LOC = "X41/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1111101001100011)
) lut_41_49 (
    .O(x41_y49),
    .I0(x39_y45),
    .I1(x38_y49),
    .I2(x39_y49),
    .I3(x39_y49)
);

(* keep, dont_touch *)
(* LOC = "X42/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010101101000010)
) lut_42_49 (
    .O(x42_y49),
    .I0(1'b0),
    .I1(x40_y49),
    .I2(x39_y47),
    .I3(x40_y49)
);

(* keep, dont_touch *)
(* LOC = "X43/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b0010011011100111)
) lut_43_49 (
    .O(x43_y49),
    .I0(1'b0),
    .I1(x40_y44),
    .I2(x40_y47),
    .I3(x41_y49)
);

(* keep, dont_touch *)
(* LOC = "X44/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000000011011111)
) lut_44_49 (
    .O(x44_y49),
    .I0(x41_y49),
    .I1(x42_y44),
    .I2(x42_y49),
    .I3(1'b0)
);

(* keep, dont_touch *)
(* LOC = "X45/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1000101100110110)
) lut_45_49 (
    .O(x45_y49),
    .I0(x43_y47),
    .I1(1'b0),
    .I2(x43_y49),
    .I3(x42_y49)
);

(* keep, dont_touch *)
(* LOC = "X46/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1011111001011011)
) lut_46_49 (
    .O(x46_y49),
    .I0(1'b0),
    .I1(x44_y49),
    .I2(x44_y49),
    .I3(x44_y44)
);

(* keep, dont_touch *)
(* LOC = "X47/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100110000101)
) lut_47_49 (
    .O(x47_y49),
    .I0(1'b0),
    .I1(x44_y49),
    .I2(1'b0),
    .I3(x44_y49)
);

(* keep, dont_touch *)
(* LOC = "X48/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b1010100000001101)
) lut_48_49 (
    .O(x48_y49),
    .I0(x45_y46),
    .I1(x46_y47),
    .I2(x45_y47),
    .I3(x45_y49)
);

(* keep, dont_touch *)
(* LOC = "X49/Y49" *)
SB_LUT4 #(
    .LUT_INIT(16'b0111110010000011)
) lut_49_49 (
    .O(x49_y49),
    .I0(1'b0),
    .I1(x47_y46),
    .I2(1'b0),
    .I3(x47_y49)
);

endmodule